brottslingar	criminals,
nederländerna	the netherlands,
andra	other,
från	from,
preussen	prussia,
buddy	buddy,
paris	paris,
tillväxten	growth,
organisation	body,
pommern	pommern,
kristendom	christianity,
ägande	ownership,
upptar	occupies,
johansson	johansson,
upplysningen	the enlightenment,enlightenment,
jack	jack,
valdes	chosen; elected,
invånare	inhabitants,
evert	everted,
stammarna	strains,
öppna	open,
chokladen	the chocolate,chocolate,
triangelns	triangle,
sydväst	southwest,
slogs	was,
sexton	sixteen,
dagens	current,
matematik	mathematics,
rollfigurer	role figure,
sovjetisk	sovietic,
parten	party,
miller	miller,
sture	sture,
sabbath	sabbath,
horn	horn,
chef	head,
alltsedan	even since,
förstaplatsen	first place,
förbättringar	improvement,
eurovision	eurovision,
indierna	indians,
bakgrunden	background,
neo	neo,
vänta	(have to) wait; expect,
unescos	unesco,
ned	bottom,
tolv	twelve,
journalist	journalist,
vampyr	vampire,
sund	healthy,
fossil	fossil,
noga	carefully,
musikalen	the musical,
flera	many,
aten	athens,
beck	beck,
parlamentariska	parliamentary,
kopplingen	the connection,
analytisk	analytical,
studeras	is studied,
sidan	page,
kategoribrittiska	category: british,
valrörelsen	the election campaign,
interstellära	interstellar,
luther	luther,
fyllde	filled,
precis	just,
dra	pull; (with)draw,
£m	million pounds,
biskop	bishop,
efterföljare	follower,
strax	just,
individerna	the individuals,
faktiskt	in fact; actually; indeed,
fördelning	distribution,
nazistiska	nazi,
slott	castle,
studioalbumet	studio album,
eftervärlden	posterity,
gävle	gävle,
betraktats	considered,
västtyskland	västttyskland,
musik	music,
giovanni	giovanni,
ljus	light,
riksväg	national highway,
ludvig	ludvig,
berlin	berlin,
lissabonfördraget	lisbon treaty,
politiker	politicians,
temperaturen	temperature,
kalksten	limestone,
kapitalistiska	capitalistic,
temperaturer	temperature,
johanssons	johansson,
ofta	usually,
utgick	was deleted,
folkmun	popular lore; popularly,
landslag	national team,
erövringen	conquest,
styrkan	strength; unit; force,
indien	india,
stommen	body,
passagerare	passengers,
genomfördes	was,
ipredlagen	ipred act,
uppmärksamhet	attention,
oavgjort	draw,
iiis	3's,
firas	celebrated,
turnera	tour,
ens	even,
gata	street,
rädd	afraid,
elektriskt	electric,
beskrev	depicted,
densitet	density,
västvärlden	western world,
gård	house,
klarar	handle,
biografen	the cinema,movie theater,
turkiet	turklet,
orden	words,
medföra	bring,
isär	apart,
lämningar	remains,
existera	exist,
liberaler	liberals,
ändra	change,
arbetslöshet	unemployment,
fifa	fifa,
vart	each,
varv	shipbuilding,
ormar	snakes,
panthera	panthera,
munnen	the mouth,
barrett	barrett,
vare	either,
organismer	organism,
besittningar	possessions,
tidpunkten	the time,
mattis	mattis,
nutida	present,
straff	penalty,
nytt	new,
wales	wales,
kanarieöarna	canary islands,
fil	file,
aborter	abortions,
avgå	resign,
startar	start,
hemlighet	secretly,
säljande	selling,
bana	web,
isen	the ice,
bank	bank,
utvecklar	development speaker,
debut	debut,
rikskansler	chancellor,
ingrid	ingrid,
laddning	charge,
café	coffeehouse,
utmed	along,
träffade	met,
voddler	voddler,
axelmakterna	the axis,
avslöjade	revealed,
daniel	daniel,
hundra	hundred,
värnplikt	military service,
standard	standard,
förmodligen	presumably,
statsöverhuvud	head of state,
inom	in,
studera	study,
ägnade	dedicated,
sannolikt	probable,
reinfeldt	reinfeldt,
sökte	searched,
professionell	professional,
starta	launch,
nätet	net,
övre	upper,
återkomst	return,
nyheten	news,
ingmar	ingmar,
starkast	strongest,
synnerligen	remarkably; particularly,
uralbergen	the ural mountains,
punkten	the point,point,
begränsar	limit,
konventionen	convention,
sång	song,
förbi	past the,
berlins	berlin's,
inget	not,
tom	tom,
uppkommit	generated,
begränsad	limited,
fördes	sea were entered,
äter	eat,
militärt	militarily,
persson	persson,
kraftverk	plant,
skildes	was seperated,
symptom	symptom,
roms	romes,
symboliserar	symbolized,symbolizes,
kontrast	contrast,
kronan	swedish krona,
sorters	kinds,
scenen	stage,
varje	each,
sheen	sheen,
regissören	director,
härkomst	provenance,
parter	sides,
minut	minute,
selassie	selassie,
folkmängden	population,
försörja	support,
värme	thermal,
stadsdelen	district,
självständiga	independent,
rak	linear,
ras	race,
fåglarna	the birds,
fasta	solid,
omvandling	transformation,
tänkt	intended,
kalendern	calender,
magnus	magnus,
lanseringen	the release,
skaffa	obtain,
sjukvård	health care,
fartyg	vessel,
muskler	muscles,
anatomi	anatomy,
närvaro	attendance,
viktig	important,
hjälpmedel	resources,
utställning	display,
bildat	formed,
fjädrar	feathers,
gallagher	gallagher,
anteckningar	notes,
thriller	thriller,
morgon	tomorrow,
dom	conviction,
freja	freja,
härstammar	derived,
sjöar	parks,
förlorar	loss,
förlorat	lost,
dos	dosage,
dop	baptismal,
singel	single,
flod	basin,
effekten	effect,
koppla	coupling,
damer	ladies,
järnvägarna	railways,
västeuropa	western europe,
bandmedlemmar	band members,
kronprins	crown prince,
vanligen	typically,
legitimitet	legitimacy,
effekter	effeckter,
rankning	rating,
sättet	way,the way,
börja	start,
teater	theater,
louise	louise,
claude	claude,
lista	list,
florens	florence,
kejsar	emperor,
breddgraden	latitude,
gärningsmannen	the offender,
helhet	entirety,
variera	vary,
holländska	dutch,
do	do,
stycke	piece; part; section,
dj	dj,
kollapsade	collapsed,
dc	d.c.,
platt	plate,
rådhus	townhouses,
watson	watson,
dy	younger,
europeisk	european,
mönster	marks,
lyssna	listening,
slags	kind,
offret	the victim,
runt	around,between,
stadskärnan	town/city,
stora	large,
existerat	existed,
bay	bay,
bad	bath,
ursäkt	apology,
fokus	focus,
release	release,
fågelarter	bird species,
kalla	cold,
ovtjarka	ovtjarka,
blev	became,
veckan	weeks,
vanlig	common,
skulle	could,
finansiella	financial,
treenigheten	the trinity,trinity,
historiens	historys,
franske	french,
arlanda	arlanda,
dittills	thus far,
ockuperat	occupied,
nuförtiden	nowadays,
djuret	the animal,
hedersdoktor	honorary doctor,
fornnordiska	old nordic,
inledningsvis	in the beginning,
månarna	moons,
sundsvalls	sundsvall,
sista	last,
finger	finder,
skrift	book,
sorts	variety,
rollen	the role,
ställning	position,
lanserades	launched,
maniska	manic,
tillämpas	applied,
muhammed	muhammed,
vinden	the wind,
fördragen	treaties,
nederlag	defeat,
svensk	swedish,
gatan	the street,
aktuell	current,
lösningsmedel	solvent,
folkmordet	genocide,
begränsade	limiting,
fångar	prisoners,
tillfälle	time,
solljus	sunlight,
varmt	hot,
basis	basis,
blodkroppar	corpuscle,
varma	hot,
socialistiska	socialistic,
patienter	patients,
life	life,
äventyr	adventure,
snittet	average,
förslag	proposal,
igång	start,
modernare	more modern,
attacker	attacks,
provinser	provinces,
chile	chile,
övergripande	overall,general,
mindre	less,
vagn	wagon,
parterna	parties,
drömmar	dreams,
invasionen	invasion,
uttryck	expression,
blåvitt	bluewhite,
grundar	bases,
kolonin	colony,
nationer	nations,
ip	ip,
förföljelser	persecution,
burundi	burundi,
dokument	files,
sommar	summer,
madonna	madonna,
nationen	the nation,
vanföreställningar	delusions,
följt	followed,
serbisk	serbian,
vänstern	left party,
vrida	turning,
kommunistpartiets	the communist party,
ernman	ernman,
gräns	limit,border,
därmed	therefore,
makt	power,
pekar	pointer,pointing,
erhållit	acquired,
hann	did,
materiell	material,
skog	forest,
hand	hand,
värde	value,
föras	taken to,
återvände	returning,
yngste	youngest,
nedan	below,
charlie	charlie,
sydamerika	south america,
glädje	joy,
rör	touch, move(-s),
centraleuropa	central europe,
mamma	mother,
monaco	monaco,
spelat	played,
grannländer	neighboring lander,
koloniseringen	the colonization,
capitol	capitol,
kraftigt	heavily,
kongressen	congress,
gods	goods,
körs	being driven,
birmingham	birmingham,
utföras	performed,
goda	good,
enades	agreed,
använt	used,
värnpliktiga	inductees,
vetenskapsmän	scientist,
julen	christmas,
eld	fire,
muhammeds	mohammed's,
huvud	main,
rätta	correct,
regionerna	regions,
född	born,
förbättra	improve,
enlighet	according,
rättegång	trial,
särdrag	feature,
svensson	svensson,
samarbete	collaboration,
föds	born,
engelskans	english,
världsdel	continent,
uppmärksammade	noticed,
hepatit	heptatitis,
sjöfarten	shipping,
läkemedelsverket	medical products agency,
årlig	yearly,
sedlar	bills,
modersmål	native language,
territorierna	territories,
studion	the studio,
gifter	toxins,
juryns	the jury's,
lagstiftningen	law-making,
vattnet	water,
hanhon	male-female,
people	people,
ansluta	join,
dead	dead,
jennifer	jennifer,
uppmärksammades	attention,
finsk	finnish,
besökt	visited,
tappar	drop,
användare	users,
princip	principle,
totala	total,
filmatiserats	been filmed,
benämns	designated,
monoteism	monotheism,
neptunus	neptunes,
angrepp	attack,
män	men,
bolt	bolt,
härstamma	stem,
annat	other; another,
därutöver	in addition,
maskiner	machines,
omgången	round,
montana	montana,
grenen	branch,
stjärna	star,
romantiska	romantic,
français	francais,
döpte	baptized,
transkription	transcription,
samer	sami,
jens	jens,
menade	meant,
psykiskt	psychic,
oförmåga	failure,
omger	surrounding,
artikeln	the article,
hantera	handle,
nova	nova,
sicilien	sicily,
jane	jane,
etablerat	established,
wittenberg	wittenberg,
form	form,
norrlands	norrland,
förhållandet	the ratio,
sagan	story,
förhållanden	relationships,
berg	mountain(-s),
verde	verde,
byggda	constructed,
finns	exist,
byggde	built,
inträffat	occurred,
gymnasiet	high school,
spelade	played,
säkerhet	safety; security,
flickvän	girlfriend,
åriga	year,
båten	boat,
beteckningen	the label,
moderna	modern,
trio	trio,
tesla	tesla,
efter	after,
handelspartner	trading partner,
tosh	tosh,
modernt	modern,
hamn	harbour,
kambodja	cambodians,
ericsson	ericsson,
förbud	prohibiting,
liberalism	liberalism,
tätorten	conurbation,
bord	table,
janukovytj	janukovytj,
dotter	daughter,
protester	protests,
arkitekter	architects,
oscar	oscar,
betalt	charge,
olja	oil,
football	football,
korrekt	proper,
jamaicanska	jamaican,
sätta	insert,
tottenham	tottenham,
katekes	catechism,
regleras	controlled,
laddade	charged,
holm	holm,
uefa	uefa,
kategorifödda	category born,
vietnam	vietnam,
rätten	right,the court,
expandera	expand,
cellens	the cell's,
skatt	tax,
funktionerna	the functions,
rob	rob,
tenderar	tend,
datum	date,
spår	track,
behöver	need,
koreanska	korean,
lider	suffers,
afrikaner	africans,
behåller	keeps,
rådet	council,
igelkott	hedgehog,
marissa	marissa,
uppdelning	division,
petersburg	petersburg,
framställa	the installation,
händelserna	events,
vladimir	vladimir,
choice	choice,
framställs	is depicted,prepared,
vegas	vegas,
skillnaderna	differences,
kusterna	coasts,
enskilt	individually,
salvador	salvador,
fackföreningar	unions,
hawaii	hawaii,
nedsatt	reduced,
hisingen	hisingen,
olyckor	accidents,
lever	liver,
säte	sate,
villa	house,
reklamen	advertising,
mån	mon,
svartån	svartån (black stream),
stimulera	stimulate,
köp	purchase,
ingick	were included,
agnosticism	agnosticism,
miniatyr	miniature,
axel	axel,
avsluta	exit,
katter	cats,
högkvarter	headquarters,head quarter,
lärde	learned,
påstår	states,claims,
avsaknad	absence,
utifrån	from,
oerhört	extremely,
spektrumet	spectrum,
huvudsakliga	main,
binder	tie,
införts	introduced,
vägg	wall,
franklin	franklin,
ankomst	arrival,
experimenterade	experimented,
bob	bob,
rafael	rafael,
diagnosen	diagnosis,
hotell	hotel,
spridit	spread,
presenterade	presented,
religionsfrihet	freedom of religion,
presenterar	present,
franco	franco,
äktenskapet	marriage,
utropades	was proclaimed,
samfundet	the communion,
samlar	salmar,
samlas	together,
vuxna	adult,
haft	had,
motsvarar	comparable,
positivt	positive,
kurder	kurds,
australian	australian,
filmer	movies,
avsattes	deposited,
flyttat	moved,
ögon	eyes,
rivalitet	rivalry,
relationerna	relations,
ställe	stalle,
hål	hole,hal,
årets	year,
kolonialismen	colonialism,
grönt	green,
tokyo	tokyo,
julius	julius,
rådgivare	advisor,
soul	soul,
allvarlig	serious,
präglade	characterized,
can	can,
generell	general,
karibiska	caribbean,
påvisa	detection,
bönorna	bean,beans,
crazy	crazy,
locka	attract,
inkluderade	included,
dennis	dennis,
kunglig	royal,
genomgått	passed,
pink	piddle,
speglar	mirror,
milda	mild,
pojke	boy,
varor	products,
till	to,
andlig	spiritual,
regeln	rule,
storleken	size,
nye	new,
kopplingar	connections,
simpson	simpson,
riktlinjer	guidelines,
löpande	conveyor (belt),
svart	black,
läkare	doctor,
upphört	end,
studenterna	the students,
natural	natural,
bergarter	rocks,
johnson	johnson,
marknad	market,
sådana	such,
romarna	the roman,
sv	south west,
tala	speak,
väntat	expected,
romantiken	romanticism,
nixon	nixon,
se	see,
väntar	expect,
resulterar	results,
komplicerad	complicated,
kong	(hong) kong,
antingen	presumably,
iberiska	iberian,
fasen	phase,
lyrik	poetry,
ingvar	ingvar,
wallace	wallace,
utsätts	exposed,
autonomi	autonomy,
äkta	married,
policy	policy,
marleys	marley's,marley,
passar	suitable,
hergé	herge,
änden	spirit,
äldste	eldest,
varav	which,
halv	half,
lejon	lion,
lagliga	legal,
spetshundar	sets dogs,
musiker	musicians,
hotar	threatens,
lockar	attracts,curls,
opera	operator,
futharkens	futhark,
stockholm	stocholm,
dominerar	dominate,
januari	january,
föremål	object,
sägs	said (to be),
födelsedag	birthday,
en	a,
greker	greeks,
valuta	exchange,
eg	ec,
förstöra	destroy,
stål	rate,
ex	eg,
eu	eu,
resultera	result,
saudiarabien	saudi arabia,
kött	cones,
åsikt	opinion,
avrättningar	execution,
årliga	annual,
riktiga	real,
bränder	fires,
brändes	burnt,
republika	republic,
bla	blah,
garantera	guarantee,
vård	nursing,
våra	our,
sålde	sells drinks,
genetisk	genetic,
juldagen	christmas day,
väster	west,
vårt	each,
dubbla	double,
california	california,
marino	marino,
brooke	brooke,
byte	change of,
nått	reached,
arbetet	work,
näring	nutrition,
sven	sven,
flandern	flanders,
massiva	massive,
artisten	the artist,
gordon	gordon,
stängdes	closed,
allmänheten	public,
någonsin	ever,
egentligen	really,
skådespelerska	actress,
satte	put together,
grupperna	groups,
fötterna	the feet,
open	open,
bergqvist	bergqvist,
skjuten	shot,
bahamas	bahamas,
skådespelarna	actors,
alfred	alfred,
grundämnen	elements,
texas	texas,
sjö	naval,
svenske	swedish,
williams	williams,
animerade	animated,
vilka	which,
användandet	use,
spelningar	gigs,
montenegro	montenegro,
alan	alan,
utrustning	equipment,
svenskarna	the swedes,
delats	divided,been awarded,
hundar	dogs,
nathan	nathan,
balans	balance,
sidorna	pages,
fiender	enemies,
ändrades	changed,
lugn	calm,
hjärtat	heart,
inträde	entry,
afrikanska	afrikanska,
tiotusentals	tens of thousands,
stadsdelar	districts,neighborhoods,
statsminister	prime minister,
kometer	comets,
faktor	factor,
formerna	forms,
grundas	based,
anger	indicates,
tänder	teeth,
hjälp	help,
övriga	other,others,
takt	rate,
förälskad	in love,
förste	chief,
fortsatta	continued,
skulptur	sculpture,
centralbanken	centralbank,
fysikaliska	physical,
potential	potential,
magnetiska	magnetic,
periodvis	periodically,
sekreterare	secretary,
tränare	coach,
successivt	progressively,
isolerad	isolation,
religionen	the religion,
förvaltning	administration,
rådets	council,
queens	queen,
över	over,
driva	run,
täckt	covered,
öppet	open,
lisbet	lisbet,
grammatik	grammar,
människan	the human,
stövare	hound,
orsaka	cause,
förfäder	ancestors,
engagemang	commitment,
axl	axl,
doktor	doctor,
nazisternas	nazi,
marocko	morocco,
tros	believed,
dahléns	dahlén's,
berättelsen	story,
guld	gold,
adolf	adolf,
himmel	heaven,
stärkte	strengthened,
ovanligt	unusual,
våld	force,
dagbok	diary,
mörk	dark,
ovanliga	rare,
analys	analysis,
depressioner	depression,
ges	given,
ger	gives,
aktiviteten	activity,
tränaren	the coach,
ambitioner	ambitions,
folkomröstning	referendum,
katla	katla (fictive dragon in the classic "bröderna lejonhjärta"),
murray	murray,
ledaren	leader,
forsberg	forsberg,
manager	manager,
försörjning	sustention,
ländernas	countries',
östblocket	the eastern bloc,
dramat	the drama,
råd	council,
roger	roger,
ljudet	the sound,
monark	monarch,
tolfte	twelth,
förmån	advantage; in favor of; benefit,
minnen	memories,
sämre	samre,
beethoven	beethoven,
drogmissbruk	drug abuse, substance abuse, drug addiction,
behovet	the need,
inspelningen	recording,
sean	sean,
slöt	joined (in peace),closed,
stanley	stanley,
minnet	memory,
menar	mean,
menas	means,
enhetlig	single,
freden	peace,
visades	showed,
federal	federal,
begränsningar	limits,
kontrakt	agreement,
kilometer	kilometers,
gaga	gaga,
människas	human,
sträcka	distance,
översättning	translation,
intresserad	interested,
ordspråk	proverbs,
hämtat	collected,
fynd	finding; finds,
antagligen	ligands presumably,
verket	board,
konstnärer	artists,
tum	inches,
comeback	comeback,
ja	yes,
värdet	the value,
vojvodina	vojvodina,
chelsea	chelsea,
ordagrant	literal,
tour	tour,
ås	ridge,
araber	arabs,
placeras	placed,
flyktingar	refugees,
pakistan	pakistan,
utnyttja	use,
cancer	cancer,
regler	rules,
syntes	synthesis,
signaler	signals,
hävda	asserting,
skånska	scanian,
sättas	turn,
överföra	transmit,
bildats	had formed,
förekomsten	presence,
luft	air,
folket	the people,
invaderade	invaded,
formen	the form,
observera	note,
skriven	written,
cobain	cobain,
elvis	elvis,
tjänster	services,
konservativa	conservative,
meningen	sense,
champions	champions,
ytan	the area,
skriver	write,
användes	was used,
bilderna	the pictures,
landskapen	the landscapes,
influenser	influences,
ansikte	face,
föregångaren	predecessor,
förlängning	overtime; extension; prolongation,
bevis	certificate,
författarskap	the writer,
pippi	pippi,
sahara	sahara,
teoretiker	theorists,
knyta	tie,
sammanfaller	coinciding,
beteckna	denote the,
ohälsa	disorders,
upplagor	issues,
långt	far,
orsakade	caused,
same	lapp,
talmannen	speaker of the riksdag,
ärftliga	genetic,
kromosom	chromosome,
träffar	hits,
samt	also,
hjärta	heart,
running	running,
linjerna	routes,
speciellt	particularly,
teknisk	technical,
lösningar	solutions,
pennsylvania	pennsylvania,
avser	regards,
värld	world,
identifiera	identification,
gudomliga	divine,
lyckan	the happiness,
berättelse	story,'s re,
koncentration	concentration,
byggnad	building,
resa	travel,
libyen	libya,
grannländerna	neighbors,
transeuropeiska	transeuropean,
programledare	host,
instrument	intrument,
spänningar	tensions,
bestämde	chose,
motverka	prevent,
lade	seized,
schwarzenegger	schwarzenegger,
underarten	subspecies,
vampyren	the vampire,
stund	while,
östergötland	Östergötland,
snart	soon,
vinkel	angle,
vampyrer	vampires,
baltiska	baltic,
skilda	separate,
patrick	patrick,
bröllop	wedding,
urval	selection,
mänsklig	human,
verksamheten	the work,activity,
lågt	low,
närheten	the vicinity,
verksamheter	activity,
strindberg	strindberg,
tiders	times,
jordbruket	the agriculture,
slår	states,
användbara	useful,
exil	exile,
cannabis	cannabis,
föra	pre,
legat	formed,
ända	up,
demokratisk	democratic,
bestämd	fixed,
willy	willy,
sätts	turned (on),
olof	olof,
nivån	level,
skär	skerry,
tyska	german,
edwall	edwall,
spelet	the game,
island	icelandic,
populationer	populations,
europeiskt	european,
torget	square,
organisationer	organizations,
upplevelser	experiences,
lands	on land,
säkerhetsrådet	security,
ansträngningar	effort,
partiet	the party,
kapten	captain,
grupperingar	groupings,
tolkning	interpretation,
burton	burton,
befinna	be,
gravid	pregnant,
satsade	bet,
klassisk	classic,
philadelphia	philadelphia,
evangeliska	evangelical,
hel	full,
hamnen	the harbour,
hänger	hanger,
gånger	times,
complete	complete,
inletts	started,
bevaras	are protected,
existerande	current,
bevarad	preserved,
gången	time,
rush	rush,
traditionerna	traditions,
expeditionen	expedition,
ingredienser	ingredient,
koenigsegg	koenigsegg,
vinkeln	angle,
miguel	miguel,
exemplar	copies,
ständig	constant,
manuel	manuel,
verkliga	fair,
regimer	regimes,
humanismen	humanism,
kostar	costs,
taylor	taylor,
ad	ad,
molekyler	molecules,
västmakterna	western powers,
bronsåldern	the bronze age,
tjorven	tjorven,
palats	palace,
väckte	aroused,
film	film,
offside	offside,
genrer	genres,
vanliga	regular,
omgivande	surrounding,
stannade	stayed,
svåra	answering,
bredare	broad,
värmlands	värmlands,
kvarstod	remained,
erövring	conquest,
henriks	henry,
vinnaren	winner,
bandmedlemmarna	band members,
symtomen	the symptoms,
villkor	conditions,
tjänare	servant,
kommunen	municipality,
kommuner	local,
århundradena	centuries,
färdas	travels,
medicinskt	medical,
snabbaste	rapid,
vila	rest,
ale	ale,
milt	mild,
vill	to,
års	years,
loppet	bore,
ingripande	negative,
zink	zinc,
ron	ron,
romanen	novel,
irak	iraq,
nederbörd	precipitation,
ögonen	eyes,
to	to,
romaner	novels,
nord	north,
cykeln	there are two meanings in the context - cycle and bicycle,
fortsatt	further,
ta	to,
ghana	ghana,
seriens	series,
ansluter	connects,
handlade	was,
fall	where,
johans	johan's,
utländsk	foreign,
uefacupen	uefa europa league,
mild	soft,
sand	sand,
siffrorna	the numbers,
sann	true,
lisa	lisa,
ockuperades	occupied,
skiva	disc,
massor	tons,
kritiserats	critized,
orgasm	orgasm,
givaren	dealer,
intressant	of interest,
höjd	height,
richard	richard,
sun	sun,
vaginalt	vaginal,
version	version,
bernhard	bernhard,
sur	sour,
sattes	was added,
islams	islams,
inblandad	mixed,
guns	guns,
lärare	teacher,
långhårig	long-haired,
fäste	bracket,attachment,
christian	christian,
dottern	the daughter,
vald	elected,
simon	simon,
medarbetare	employees,
traditionella	traditional,
stulna	stolen,
minst	at least,
boxning	boxing,
känsliga	susceptible,
social	social,
alice	alice,
globen	lobe,
vid	at,in,
snus	snuff,
nazityskland	nazi germany,
uppkomst	origin,
grunda	base,
stöd	support,
juridiskt	juridical,
varianterna	variants,
avsedd	intended,
spelaren	the player,
socialdemokraterna	members of the social democracy,
biskopen	bishop,
rösterna	votes,
tillät	allowed,
spelades	filmed,
representerar	represents,
rhen	rhine,
massan	mass,
mord	murder,
ragnar	ragnar,
utökat	expanded,
alltid	always,
latinamerikanska	latin american,
människa	man,
brist	non,
uppskattas	estimated,
räknas	counted,
gogh	gogh,
glad	happy,
berätta	tell,
medelklassen	middle class,
science	science,
mördad	murdered,
företeelser	phenomena,
sociala	social,
den	it,
befintliga	current,
samtliga	all,
history	history,
skadliga	deleterious,
varelse	creature,
huvudstaden	capital,
mellersta	middle,
feministiska	feminist,
betoning	stress,
spansk	spanish,
medförde	led,
sträng	strang,
stil	type,
sålts	sold,
gälla	valid,
rapport	report,
uppnått	met,
uttrycka	express,
begränsa	limit,
samarbetet	cooperation,
hoppade	jumped,
fortsättning	further accession,
torde	should,
försök	expirements,
referens	reference,
lanka	(sri) lanka,
köpte	bought,
vattenkraft	water power,
bildade	formed,
pucken	the puck,
kognitiv	cognitive,
segrar	wins,
kategoriorter	category visited,
rockgrupper	rock groups,
greklands	greek country,
komplexa	complex,
nämnts	mentioned,
bernadotte	bernadotte,
avvisade	rejected,
blommor	flowers,
gudarnas	gods,
göra	do,
mörkt	dark,
färöarna	the faroe islands,
länge	long,
mörka	dark,
vietnamkriget	vietnam war,
islam	islam,
rika	rich,
protestanter	protestants,
caesars	caesars,
edmund	edmund,
stephen	stephen,
epok	epoch,
argentina	argentina,
jämte	together with,
good	good,
otto	otto,
musikalisk	musical,
bytte	changed it's,
kärna	quarks,
säkerhetsråd	security council,
dyrt	a high price,expensive,
grekisk	greek,
närmare	further,
landborgen	the ridge,
marcus	marcus,
exemplet	example,
intåg	entry,
kungarna	kings,
slidan	the vagina,
skrivit	written,
lägre	lower,
härrör	derived,
enstaka	occasional,
michael	michael,
energy	energy,
doser	dose,
aldrig	never,
energi	energy,
kretsen	the order,
sexuella	sexual,
sanningen	truth,the truth,
nationens	the nation's,
oftast	usually,
infrastrukturen	the infrastructure,
research	research,
ölet	the beer,
uppstått	arised,
fullständig	complete,
kopplat	coupled,
sparken	park,
stöder	supports,
känna	known,
strömning	strom accession,
vikingar	vikings,
ålands	the Åland island's,
eventuellt	eventually,
delningen	division,
viken	gulf,
bära	carry,
polisen	the police,
faller	fall,
målningar	paintings,
utöver	addition,
ytterligare	further,additional,
sändes	sent,
elden	the fire,
riksföreståndare	regent,
spekulationer	speculations,
fabriker	factories,
bland	inter,
kol	coal; charcoal,
avel	breeding,
parlamentsvalet	parliamentary elections,
sår	wound,
brasiliens	brazil's,
förhindrar	prevents,
familjerna	families,
brittiska	british,
traditionen	the tradition,
brittiske	british,
gränser	borders,
åkte	went,
kardinal	cardinal,
modet	the fashion,
järnvägar	rail,
hotet	the threath,
fattigaste	poorest,
zeppelin	zeppelin,
influerad	influenced,
matteusevangeliet	book of matthew,
humanistiska	humanistic,
king	king,
fattiga	poor,
direkt	direct,
organiserat	structured,
nöd	distress,emergency,
knapp	scarce,
andersson	andersson,
värden	values,
personens	the persons,
haddock	haddock,
hellström	hellström,
stiftelsen	foundation,
följder	impact,
äga	own,
kusin	cousin,
gjort	created,
karl	karl,
vädret	the weather,
visats	demonstrated,
publicerad	published,
kongokinshasa	kong kinshasa,
genast	immediately,
varianter	diversities,
avseenden	regard,
victor	victor,
mexiko	mexico,
lettland	latvia,
hotel	hotel,
dagliga	daily,
säsongens	season,
naturvetenskapliga	scientific,
bistånd	aid,assistance,
dagligt	daily,
utbrott	outbreaks,
part	party,
klädd	coated,
microsoft	microsoft,
statsskick	government,
thomas	thomas,
tjugo	twenty,
lön	salary,
karaktär	character,
ursprungliga	original,
kolonialism	colonialism,
antagit	adopted,
richmond	richmond,
konto	account,
svenskans	the swedish language,swedish language,
befolkningstätheten	population density,state of the population,
canaria	canaria,
indian	indian,
rädsla	fear,
ikon	icon,
världens	the worlds,
lennon	lennon,
igelkottar	hedgehogs,
jämfört	compared to last,
ingå	include,be included in,
beyoncé	beyoncè,
beslutar	decides,
vänskap	friendship,
tekniken	techinque,
jobbade	worked,
händer	happens,
förklarar	explains,
restauranger	restaurants,
stadsparken	city park,
skapelse	creation,
vincent	vincent,
river	tear,
etiopien	ethiopia,
ser	see,
maurice	maurice,
suveränitet	sovereignty,
vind	wind,
tidigare	earlier,
are	are,
järnväg	rail,
sen	then,
stjäla	steal,
nations	nation,
institutet	institute,
barn	child,
guden	god,
chefen	commendant; commander,
bortsett	except,
planerar	plan,
lösa	solve,
fission	fission,
löst	dissolved,
europe	europe,
läns	county,county's,
romarriket	the roman empire,
latin	latin,
iron	iron,
framfört	presented,
allvar	serious,
intäkter	incomes,
rösten	rust,
uppkom	arose,
skivorna	plates,
produkter	products,
statligt	governmental,
tiderna	the times,
uppfattning	view,
roman	novel,
restaurang	restaurant,
använda	using,
bott	lived,
globala	global,
omkom	perished,
kroatiens	croatia's,
uppfylla	fulfill,
andas	breathes,
således	hence,
scientologikyrkan	the church of scientology,
immunförsvar	immune defense,
stärktes	strengthened,
church	church,
natt	night,
skydd	protection,
hypoteser	hypotheses,
ps	p.s,
minskade	minimum period,
våningar	floors,storeys,
oändligt	infinitely,
laos	laos,
gestalt	character,
beskrevs	described,
isolerade	isolated,
gav	gave,
togs	taken,
anthony	anthony,
livet	life,
uppleva	experience,
kalmar	kalmar,
bild	picture,
konflikter	conflict,
läses	read,
brottslighet	crime,
arenan	arena,
ris	rice,
titanic	titanic,
rik	rish,rich,
korruptionsindex	corruption perceptions index,
hovet	court,
barney	barney,
borgerliga	conservative,
sjuk	ill,disease,
omvandlas	converted,
skalet	the shell,
högste	highest,
förföljelse	persecution,
dödad	killed,
omgivning	surroundings,ambient,
tyder	indicates,
arméer	armies,
luxemburg	luxemburg,
skeppet	the ship,
byar	villages,
uppbyggd	structered,
debatter	debates,
republiker	republics,
uppbyggt	structured,
debatten	the debate,
vargar	wolves,
euro	euro,
älska	love,
kurdisk	kurdish,
normala	normal,
albanien	albania,
italiensk	italian,
skildringar	description,
normalt	normally,normal,
person	person,
edge	edge,
johan	johan,
följande	the following,
ande	of,
njurarna	kidney,
senaste	last,
alternativt	alternatively,
skal	shell,skin,
påverkade	affected,
remmer	remmer,
kallblod	draught horse,
taiwan	taiwan,
tropisk	tropical,
sektion	section,
namnet	the name,
sparta	sparta,
fascistiska	fascist,
minoriteten	minority,
nordväst	north west,
jönssonligan	jönssonligan,
namnen	the names,
pornografi	pornography,
marco	marco,
teknik	technic,
kulturen	the culture,
inkomsterna	revenue,
baserade	based,
rastafarianerna	the rastafarian,
bit	piece,
rené	rené,
releasedatum	release date,
dylikt	such,
banbrytande	groundbreaking,
gandhis	gandhi,
terminologi	terminology,
informationen	the information,
hittat	found,
minskning	reduction,decrease,
begärde	called,
norrut	north,
tål	stand,
sjöfart	maritime,
betraktar	sees,
jordbävningar	earthquakes,
utvecklades	developed,
läste	read,
ungefär	approx.; approximately,
höjden	height,
sammanhängande	connective,
måste	must,
statyn	the statue,
per	per,
kejsarens	emperors,
be	be,
bl	short of "bland" - in the context: bl. a (bland annat) = among others,
palmes	palme's,
ställningen	position,
anklagades	accused,
santa	santa,
kostnaderna	costs,
russell	russell,
bosättningar	settlements,
gemenskaperna	communities,
tätt	tight,
britannica	britannica,
vägarna	paths,
fungerande	effective,
oktoberrevolutionen	the october revolution,
clinton	clinton,
anföll	attacked,
syret	oxygen,
hemingway	hemingway,
styrelse	board,
kravet	requirement,
ön	the island,
steven	steven,
reglerna	rules,
ordnar	decorations,
hållet	cohesive,
paret	parathyroid,
befolkningens	population's,
överst	top,
dröja	wait,
ligga	lie,
visar	shows,
dalar	valleys,
samerna	sami,
turkiska	turkish,
rasade	collapsed,
regionen	region,
begreppen	the terms,
jaga	course,
sköter	handle,
serie	series,
konsul	consulting,
begreppet	the term,
samlag	intercourse,
cia	cia,
anklagelser	allegations,
mångfald	variety,
eviga	eternal,
styrande	rulers,
ur	from,
källa	source,
erövrades	(was) conquered,
trafikerade	frequent,
planer	plans,
förbjöds	banned,
reggaen	reggae,
jordbävningen	earthquake,
tropiskt	tropical,
dog	died,
skandinavien	scandinavia,
personlighetsstörning	personality disorder,
eller	or,
edwards	edwards,
sjunde	seventh,
hanen	the cock,
musikens	music,
matematiker	mathematician,
berättas	is told,
skyddas	skyas,
individuella	individual,
feodala	feudal,
besegra	defeat,
dominerades	was dominated,
inkomstkälla	source of income,
djurgårdens	djurgården's,
medina	medina,
regissör	director,
nådde	reached,
jagar	hunting,
slås	slas,
modernismen	modernism,
judisk	jewish,
delta	participate,
nasa	nasa,
regionalt	regional,
folkliga	popular,
tungt	heavy,
dvs	d.v.s.,
indiska	indian,
sitta	sit,
företeelse	feature,
sigmund	sigmund,
låter	let,
lilla	small,
hindra	prevent,
hamnar	ports,
hamnat	got,got in to,
konsten	art,
monoteistiska	monotheistic,
sent	late,
luleå	luleå,
kategoritvseriestarter	category television series starts,
märken	brands,
presidentens	the president's,
kedjan	the chain,
kommunistiska	communist,
rinner	flow,
utgjordes	make up,
vägrade	refused,
befälhavare	commander,
svts	svts,
tillhörande	associated,
tro	believing,
påverka	impact,
byggt	built,
tre	three,
utanför	outside,
leonardo	leonardo,
socialdemokratiska	social democratic,
joey	joey,
storhetstid	heyday,
bolsjevikerna	bolsevikema,
förlust	loss,
sändas	sent,
överhöghet	suzeranity,
geologiska	geological,
skadan	the hit,
direkta	direct,
ställde	asked,
årtionden	decades,
börjat	begun,
västlig	western,
konstant	constant,
depression	depression,
kinas	kinase,
hölls	was,
går	is,
chicago	chicago,
bjöd	offered,invited,
gradvis	progressively,
praktiken	effectively,practically,
indiens	indias,
tillkomst	established,
krig	war,
ledande	conductive,
utrikespolitiken	the foreign policy,
journal	jurnal,
offentlig	public,
lee	lee,
extremt	extreme,
eminem	eminem,
åtgärder	measures,
uppgick	total,
ryska	russian,
händelser	handelsar,
innebandy	floorball,
talang	talent,
störning	noise,high accession,
medeltid	medieval,
metro	metro,
tegel	brick,
krönika	chronicle,
västerut	westward; west,
chans	chances,
plattan	the plate,
opinion	opinion,
existens	existence,
talare	speakers,
hennes	her,
nås	reached,
distriktet	district,
betraktas	considered,
medlemsstater	member,member-state,
varpå	thereafter,
kinesisk	chinese,
personen	person,the person,
tas	is taken,
hemlig	secret,
utdöda	extinct,
klaviatur	keyboard,
stärka	strengthen; bolster,
nytta	good,
orkester	orchestra,
inlandet	inland,
författning	constitution,
ytterst	highly,
öppnat	opened,
andliga	spiritual,
invigningen	inauguration,
införande	introduction,
hindrade	prevented,
ansvaret	the responsiblity,
fungerar	works,
gabriel	gabriel,
advokat	bar,
avseende	regard,
beskrivs	described,
kenny	kenny,
monica	monica,
process	process,
ledamöterna	the commissioners,
hilton	hilton,
tryckta	printed,
beslöt	resolved,
saken	the matter,
hercegovina	herzegovina,
fördelningen	distribution,
föregående	preceeding; previous,
gitarr	guitarr,
romantikens	romanticism,
saknade	lacked,
tågen	the trains,
internationella	international,
undantaget	except,
revs	was demolished,
böckerna	books,
dramaten	dramaten,
gunwer	gunwer,
väpnad	armed,
trycktes	printed,
kontroversiellt	controversial,
herrlandskamper	men's international contests,
dödlig	lethal,
fart	off,
tack	thanks,
klan	clan,
gammal	old,
terrier	terriers,terrier,
diskuterades	discussed,
strategiska	strategic,
väckt	woken,
dryck	beverage,
slutsatsen	the conclusion,
registrerade	data,
mekka	mecca,
obelix	obelix,
olyckan	the accident,
offentliga	public,
riktningen	direction,
blandas	mixed,
spotify	spotify,
belopp	amounts,
frivilliga	volunteers,
glenn	glenn,
byn	village,
spanjorerna	spaniards,
tecknet	the sign,
föreställer	depicts,
uppdelad	split,
uppmärksammat	attention,noticed,
filosofiska	philosophical,
verkligen	the reality,
dag	dag,
utfärdade	issued,
bryter	breaks,
avslöjar	reveals,
tillkommit	been,
försämrades	decreased,
periodiska	periodic,
satelliter	satellite,
bas	base,
sönder	probes,
exempelvis	e.g.,
delat	divided,
vidta	take,
australiska	australian,
juridisk	legal,
krita	chalk,
företrädare	representatives,
smallwood	small wood,
fördrevs	ford described,
intresset	interests,
uppfattas	be perceived,
etymologi	etymology,
borderline	borderline,
minskad	reduced,
kärnan	core,
hantverkare	craftsman,
fiktiva	fictitious,
huvudstad	capital city,
bål	torso,
nobelpristagare	nobel laureate (-s); nobel prize winner (-s),
plural	plural,
upphörde	expired,
hjälpt	helped,
höra	hear,
uppe	top,up,
förstod	understood,
arbetare	workers,
förändra	change; alter; replace,
kortare	shorter,
florida	florida,
blanda	mix,
adrian	adrian,
tigrar	tigers,
ifrån	off,
kräva	demand,
stämmer	(if it's) true,is true,
pga	because of (short of "på grund av"),
användningsområden	possible use,
önskemål	desire,
regenter	monarchs,
skyddade	protected,
därav	thereof,
nätverk	network,
studerade	studied,
nationalistiska	nationalist,
leder	leads,lead,
spaniens	spain's,
fågelhundar	bird dogs,
omfattning	extent,
mao	mao,
rösträtt	right to vote,
kuben	the cube,
havet	sea,
belgiska	belgian,
hasch	hashish,
sjögren	sjögren,
konservativ	conservative,
släkten	genera,
bevarats	preserved,
franska	french,
domaren	the judge,
inne	inside,
light	light,
premiär	premiere,
bet	bit,
samverkan	co,
jonatan	jonathan,
stöds	stood,
tids	time,
operativsystem	operative systems,
kvinnans	female,
jämförelsevis	comparative,
flyttar	move,
vända	turn,
farligt	dangerous,
byggas	prevented,
följs	followed,
uppfann	invented,
min	my,
mills	mills,
filosofin	philosophy,
sinatra	sinatra,
besättningen	crew,
konstverk	artwork,
praxis	practice,
attackerna	the attacks,
centre	centre,
runorna	the runes,
röst	voice,
förblev	remained,
jorge	jorge,
dinosaurier	dinosaurs,
missionärer	missioners,
visa	see,
genomslag	impact,
resultaten	the results,
öken	desert,
upprustning	renovation,
irakkriget	iraq war,
republikanska	republican,
nordöst	northeast,
judendomen	the judaism,
synligt	visible,
skogar	forests,
viktigaste	most important,
styrka	strength,
text	text,
debatt	debate,
inhemsk	native,
fynden	finds; findings,
ugglas	ugglas,
bussar	bus,
euroområdet	euro area,
fursten	prince,
jan	jan,january,
shahen	shah,
varit	been,
beroende	depending,
partnern	partner,the partner,
skarsgård	skarsgård,
piratpartiet	pirate party,
klassiska	classic,
buddhismen	buddism,
inbördeskrig	civil war,
lägger	lies,
lucky	lucky,
inflytelserika	influential,
generalen	the general,
parlamenten	the parliament,
linje	line,
klassiskt	classic,
uppehåll	residence,
kämpade	decreased,
närstående	relatives,kindred,
tidigaste	earliest,
britterna	the brits,
fuglesang	fuglesang,
vänt	turned,
national	national,
svenska	swedish,
priset	the prize,
kronisk	chronic,
uppträdde	occurred,
svenskt	swedish,
först	first,
mestadels	most of the time,
reform	reform,
konverterade	converted,
rikare	richer,
upprättandet	establishment,
carlsson	carlsson,
avslutades	closed,
företagets	the corporation's,
ken	ken,bank,
balansen	balance,the balance,
finalen	final,
satsa	bet,
hårdare	more severely,
merry	merry,
jobba	work,
förklaringar	explanations,
jon	jon,
kedjor	chains,
hits	hits,
empathy	empathy,
allsvenskan	headlines,
påtagligt	markedly,
fåglar	birds,
framgångsrika	succesful,
april	april,
belägen	disposed,
älskar	loves,
kommendör	commander,
klasser	classes,
helsingfors	helsinki,
exakta	exact,
korruption	corruption,
dör	dies,
wall	wall,
utsågs	was appointed,
död	dead,
johann	john,
stabila	stable,
publiceras	will be published,
kings	kings,
dök	appeared,turned,
publicerat	published,
liberala	liberal,
antal	number of,
klara	clear,
hindu	hindu,
sara	sara,
månar	moons,
äldre	old,older,
slippa	avoid,
växt	plant,
strindbergs	strindberg,
antas	is required,
define	define,
mike	micke,
pontus	pontus,
dominera	dominate,
affärer	business,
stationer	stations,
spaniel	spaniel,
fortsättningen	remain,the continuation,
ätten	the dynasty,
sänts	sants,
strömningar	tendencies,
gärning	deed,
därifrån	from thence,
huvudet	head,
bråk	fraction,
officiell	official,
bruket	use,the use,
mandatperiod	term (of office),
långsamma	slow,
klassificera	classifying,classify,
platons	platon's,platos,
nordens	the scandinavian countries',
cypern	cyprus,
vd	ceo,
förlopp	pattern,developments,
demo	demo,
vm	vm,
flickor	girls,
måleri	painting,
vistelse	stay,
föreligger	is,
röra	move,
spela	play,
tupac	tupac,
huden	skin,
paulo	paulo,
buddhism	buddhism,
förebyggande	preventive,
känd	known,
terrorism	terrorism,
skickade	sent,
kustlinje	coastline,
övervägande	the predominant,
hinduismen	hinduism,
införa	introducing,
framförde	performed,
helsingborgs	helsing borg,
infört	introduced,
rätt	steering wheel,
kallar	calls,
alperna	alps,
strömmen	the stream,
banden	bands,
omgångar	cycles,
banker	banks,
agnostiker	agnostics,
hårdrocken	hard rock,
onda	evil,
kontakt	plug,
paus	pause,
singeln	singeln,
sänds	sands,
möjligheter	potential,
sofie	sofie,
förekommer	occurs,
patrik	patrik,
jarl	earl,
kampf	kampf,
hoppa	skip,
lära	get to know,
engelsk	english,
nacional	nacional,
ska	will,
framtid	future,
match	game,
psykoser	psychoses,
jesper	jesper,
motorvägen	highway,
vanligare	more common,
historia	history,
definitivt	unavoidable,
know	know,
klassificering	classification,
lincoln	lincoln,
lär	learn,
koden	the code,code,
vallhund	herder,
djupa	deep,
amazonas	amazonas,
sarajevo	sarajevo,
works	works,
uppträda	appear,
nationalpark	national park,
trotskij	trotskij,
starkaste	strongest,
förlusterna	the losses,
aktier	stock,
förenklat	simplified,
försvinna	disappear,
peter	peter,
transport	carriage,
skriftliga	written,
planering	planning,
joachim	joachim,
stieg	stieg,
behandlades	treated,
låten	song,
toppar	(that) peaks,
löser	solves,
skildrar	portrays,
knä	knees,
ledd	led,
fristående	independent,stand-alone,
internationalen	international,
svaga	faint,weak,
halvön	the peninsula,
ateism	atheism,
östberlin	east berlin,
sommarspelen	summer olympics,
usas	u.s.,
smärta	pain,
vargen	the wolf,
substantiv	noun,
freedom	freedom,
glada	happy,
bestämma	determining,
andel	share,
aspergers	aspergers,
samlats	solid,
troligen	probably,
reaktionerna	the reactions,
armar	arms,
alexanders	alexanders,
förstärka	enhance,
socken	parish,
anpassade	custom,
tränger	forces forward,
sekelskiftet	the turn of the century,
räddade	saved,
tendenser	tendencies,
mera	more,
vimmerby	vimmerby,
glukos	glucose,
observatörer	observers,
vad	what,
djävulen	the devil,
skola	school,
blå	blah,
regisserad	directed,
vacker	beautiful,
bedöms	evaluated,
förändrades	changed,
distinkt	distinctive,
påverkat	affected,
cricket	cricket,
radioaktiva	radioactive,
granne	neighbour,
neutral	neutral,
hundratal	hundred,
ersättning	pay,
hc	h.c,
ha	have,
radioaktivt	radioactive,
svält	starvation,starvations,
nöjd	content,
volvo	volvo,
allierad	allied,
tema	theme,
ovanför	over,
vänstra	left,
bitar	bit,
beatrice	beatrice,
stormakter	world powers,
heter	is named,
bosättare	settlers,
paraguay	paraguay,
utnyttjar	uses,
skilsmässa	divorce,
separerade	separated,
manlig	male,
året	all year,
sänktes	reduced,
särskilda	special,
proteinet	the protein,
ep	ep,
relationen	ratio,
fattigdomen	poverty,
åren	the years,years,
övergång	transition,
huvudstäder	capital cities,
shakespeares	shakespeare's,
tvfilm	tv-movie,
ställningar	notions,
kritik	critisism,critique; criticism,
variation	diversity,
koncentrationsläger	concentration,
färgerna	colors,
stad	city,
musikvideon	music video,
flyger	flying,
philips	philips,
vana	used,
stadens	the citys,city's,
etiken	ethics,
framför	above,
påverkar	affecting,
blogg	blog,
