vanligast	most,most usual,most common,
nordisk	norse,nordic,
uppemot	almost,up,
stammarna	tribes,strains,
arternas	the species,species,
jihad	johad,jihad,
elva	eleven,
invandrare	immigrants,immigrant,
hållas	be,be held,
albumet	album,
slå	beat,hit,
albumen	the albums,albums,
hermann	hermann,
lord	lord,
vann	won,
lyckats	succeeded,
dela	divide,dividing,
katoliker	catholics,
organisation	body,organization,
regional	regional,
upptar	occupies,
lämnades	was lefted,was,left,
portugals	portugals,portugal,
dels	and,both,partly,
skicklig	skillful,proficient,skilled; skillful,
statlig	state,government,
medelhavet	mediterranean sea,mediterranean,
andre	other,
helsingborg	helsingborg,
haber	haber,
befogenheter	authorities,powers,
triangelns	triangle,the triangle's,
urskilja	distinguish,discern,
sovjetisk	soviet,sovjetic,sovietic,
miller	miller,
sture	sture,
sammansatta	composite,composed,joined,
selassie	selassie,
ungerns	hungary,hungrarys,hungary's,
hanar	males,
upprätthåller	maintains,maintaining,
åsikten	the opinion,view,
åsikter	opinions,
breddgraden	latitude,parallel,
fossil	fossil,
koffein	caffeine,caffein,
jönsson	jönsson,johnsson,
filosofer	philosophers,philosopher,
aten	athens,
hårda	hard,
biografi	biography,
vägrar	refuses,refuse,
filosofen	the philosopher,
motståndsrörelsen	the resistance,resistance,
regnskog	rain forest,rainforest,
herr	mister,mr,
föräldrarna	the parents,parents,
valrörelsen	election campaign,
bipolär	bipolar,
kids	kids,
demokratier	democracies,
naturen	the nature,nature,
blåser	blows,blowing,
vicepresident	vice president,
robin	robin,
miljarder	billion,billions,
karin	karin,
tillverkningen	production,the production,
snö	snow,
unik	unique,
norsk	norwegian,
iis	ii's,
marino	marino,
hamas	hamas,
systematiskt	systematically,systematic,
ansluta	join,connect,
dna	dna,
sjukdomen	disease,
strikt	strict,
fuktiga	damp,damply,
betraktats	considered,been seen,(been) viewed,
music	music,
dns	dns,
fuktigt	moist,damp,humid,
gallien	gaul,
musik	music,
befolkningstillväxten	population growth,the population growth,the growth of population,
mercurys	mercury's,mercurys,
holm	holm,
politiker	politicians,politician,
slutligen	back end,finally,at last,
bulgariska	bulgarian,
temperaturen	temperature,
kalksten	limestone,
teman	themes,
temperaturer	temperature,
ofta	usually,often,
avancerad	advanced,
vännen	the friend,friend,
köpa	purchase,buy,purchasing,
befolkningsutveckling	population development,population growth,
vågen	the wave,scale,
stommen	body,frame,the foundation,
köpt	purchased,bought,
passagerare	passengers,passenger,
kapitalismen	capitalism,
want	want,
absoluta	absolute,
vänner	friendas,friends,
igelkottar	hedgehogs,
hon	she,
kallare	colder,
hov	court,
how	how,
hot	hot,
pågick	lasted,
folkmusik	folk music,
typen	model,the type,type,
fylla	fill,
inrikes	domestic,
trettioåriga	13 year olds,thirty year's (war),thirty years,
barbro	barbro,
sedd	seen,
objekt	objects,object,
turkiet	turkey,turklet,
sankt	st.,sankt,
typer	characters,types,
stormaktstiden	great power period,greatness,
grekiska	greek,
isär	ice,apart,
arbeten	works,
deutsche	deutsche,
hemlandet	the home country,the homeland,
wind	wind,
blind	blind,bank,blank,
varv	revolutions,dockyard,shipbuilding,
ormar	snakes,
vars	whose,who's,
dalí	dali,
organismen	the organism,organism,
vare	either,
varg	wolf,
organismer	organism,organisms,
vara	be,
barnet	child,
mabel	mabel,
varm	hot,warm,
publicerade	published,
besläktade	related,
nutida	present(-day); contemporary,present day,present,
wales	wales,
målade	painted,
assyriska	assyrian,
fil	master of,file,
avgå	resign,
väte	hydrogen,
hemlighet	secretly,darkness,
säljande	selling,
bestämmer	determines,decide,
hänga	hang,
närliggande	adjacent,nearby,
silver	silver,
utvecklat	developed,evolved,
utlänningar	foreigners,
utvecklar	develops,development speaker,
utvecklas	development,
terrorister	terrorists,
tingslag	leet,things type,
debut	debut,
utveckling	development,
tillgängligt	available,
utvecklad	developed,
andrew	andrew,
ingrid	ingrid,
tillgängliga	available,
uppnådde	met,achieved,
talade	spoken,spoke,
sapiens	sapiens,
lätt	easy,
serier	comics,series,
allan	allan,
utvecklandet	development,
serien	series,the series,
truman	truman,
axelmakterna	the axis,axis,
varken	neither,either,
kontrollerade	controlled,
slovenien	slovenia,slovenian,
försökt	tried,
förändringar	changes,
foundation	foundation,
debatter	debates,
nuvarande	current,
anarkister	anarchists,
metallica	metallica,
arbetsplats	work,workplace,
ägnade	dedicated,
sannolikt	probably,probable,
att	to,that,
sysselsätter	employs,
atp	atp,
okända	unknown,
malmös	malmö's,malmö,
sydost	south east,southeast,
givetvis	course,naturally,
grannlandet	neighboring,the neighbouring country,
östberg	Östberg,ostberg,
tecknade	cartoon (-s),cartoon,drew,
övre	upper,top,
ledarskap	leadership,
förespråkar	advocate,advocates,
xii	xii,
xis	the eleventh's,
master	masters,master,
vågade	dared,
ära	oar,glory,honor,
bitter	bitter,
förändringarna	changes,change,
senaten	senate,the senate,
bokstäverna	the letters,letters,
förmögenhet	fortune,wealth,
placerade	put,placed,placed (in),
nirvana	nirvana,
påverkad	influence,affected,influenced,
ahmed	ahmed,
skatter	taxes,
upphov	origin,source,rise,
tyckte	thought,found,find,
påverkan	impact,influence,
tree	tree,
upplysningstiden	enlightenment,age of enlightenment,
nations	nation,nations,
trey	trey,
varje	each,
utformningen	the layout,layout,the design,
påverkas	affected,
tretton	thirteen,
obligatorisk	obligatory,mandatory,
folkmängden	population,
försörja	support,
assistent	assistant,
kriterierna	criteria,
boston	boston,
dricker	drinking,drink,drinks,
filosofisk	philosophical,philosophic,
halva	half,
joakim	joakim,
trakten	the region,region,area,
fasta	solid,firm; set; solid; fast; fasting,
kroatien	croatia,
normalt	normally,normal,
östeuropa	eastern europe,east europe,
skaffa	get,obtain,gain,
spelningar	tour,gigs,
dikter	poems,
förhärskande	dominant,prevailing,
himlen	heaven,although the sky,
hjälpmedel	aid,resources,means agent,
bedrivs	conducted,
katalonien	catalonia,
konserthus	concert hall,concert,
victoria	victoria,
gallagher	gallagher,
medlemsstaterna	member,member states,
anteckningar	notes,
bedriva	carry,prosecute,
eftersom	while,because,
thriller	thriller,
övertog	took over,overtook,
annars	else,
singer	singer,
morgon	tomorrow,morning,
arkitektur	architecture,
öland	oland,öland,
camp	camp,
utmärkande	characteristic,distinguishing,
förlorar	loss,loses,
översatt	translated,the translation,
förlorat	lost,
producent	producer,
grovt	heavy,rough,roughly,
passerade	passed,
singel	single,
tänkte	thought,was going to,
inspelning	recording,
ungar	kids,babies,kids; offsprings; young,
representanter	represenatives,representatives,
bomb	bomb,
bandmedlemmar	band members,
diplomatiska	diplomatic,
sannolikhet	probability,
pris	price,prize,
teater	theatre; theater,theater,
louise	louis,louise,
populärkultur	popular culture,pop-culture,
buss	bus,
than	than,
övergår	surpasses,released,exceed,
rico	rico,
bush	bush,
omvända	reverse,
rice	rice,
mottog	received,
lastbilar	truck,trucks,
storbritanniens	united kingdom,uk,
tillståndet	state,condition,the state,
rättegången	trial,the trial,
årsdag	anniversary,
metoder	methods,
upprätta	establish,up,
metoden	the method,
dansk	danish,
plats	place,spot,place; position,
nathan	nathan,
lyssna	listening,listen,
begravning	funeral,
innebörd	meaning,
spänning	voltage,
hantverk	crafting,crafts,
×	x,
kallt	cold,coldly,
sköta	manage,operate,handle,
utgåvan	edition,issue,the edition,
uppgift	task,data,
framfördes	framfordes,were,
kontroll	control,
sköts	postponed; run,shot,handled,
kalla	cold,
ovtjarka	caucasian shepherd dog,
blev	became,was,
etik	ethics,
flagga	flag,
skulle	could,would,
skriva	write,
bygger	based,(is) building (on),
arlanda	arlanda,
skrivs	written,printed,
nuförtiden	nowadays,today,
hedersdoktor	honorary doctor,honorary degree,honorary doctorate,
manson	manson,
förhindra	prevent,
wikipedia	wikipedia,
upphovsrätt	rise knob,copyright,
sundsvalls	sundsvall,(city of) sundsvall's,
figur	figure,
sista	last,
siste	lattermost,last,
pirate	pirate,
ringa	call,
rollen	role,the role,
henrik	henrik,
ställning	position,
lanserades	launched,was launched,
tilldelades	awarded,
kommunikation	communication,communications,
världsturné	world tour,
roller	roles,
kloster	monastery,
tillämpar	administer,practice,administers,
tillämpas	applied,
huvudet	head,the head,
country	country,
kubas	cuba's,cuba,
följas	followed,
pitt	pitt,
edgar	edgar,
nordiska	nordic,
underlätta	ease,facilitate,
anordnas	provided,arranged,organised,
nordiskt	nordic,
genus	gender,genus,
logik	logic,
summan	sum,the sum,
igelkotten	the hedgehog,hedgehog,
folkmordet	genocide,
armén	the army,
uttal	pronunciation,pronounciation,
baháulláh	bahaullah,bahullah,
afrikanska	afrikanska,african,
fra	fra,
union	union,
avgörande	settling,decisive,essential,
fri	free,
anc	anc,
operationer	operations,
socialistiskt	socialistic,socialist,
årtionde	decade,
fru	madam,mrs.,wife,
arbetslösheten	unemployment,
verktyg	tool,tools,
barndom	childhood,
life	life,
café	cafe,coffeehouse,café,
snittet	average,the intersection,the average,
huvudstäder	capital cities,capitals,
ändrade	changed,modified,
arkiv	archives,archive,
närvarande	present (-ly),present,
dave	dave,
kometer	comets,
chile	chile,
övergripande	over arching,overall,general,
chili	chili,
parterna	parties,
intag	intake,
slutliga	evenutal,final,ultimate,
frankrikes	frances,france's,
castro	castro,
klarade	made it,passed,
organisera	organize,organizing,
kontraktet	the contract,contract,
tintin	tintin,
k	k,
åke	åke,
brister	failures,inabilities,
gärna	i'd love to,readily,
desto	the,ever,
stämma	sue,meeting,
player	player,
fascismen	the fascism,fascism,
australia	australia,
bristen	lack of,lack,
slag	kinds,type,
madonna	madonna,
tät	compact,sealed,frequent,
memorial	memorial,
serbisk	serbian,
tillhandahåller	provides,
vrida	twist,turn,turning,
foton	images,photos,
omkring	surrounding,about,around,
agnetha	agnetha,
european	european,
materiell	material,
klimatet	environment,climate,the climate,
josef	joseph,josef,
topp	top,
värde	value,
emi	emi,
tunn	thin,
föras	be,be brought,taken to,
synder	sins,
tung	heavy,
obligatoriskt	obligatory,mandatory,
finska	finnish,
lucas	lucas,
kampanj	campaign,
centraleuropa	central europe,
gudinnan	goddess,the godess,
grundlag	constitution,
misslyckade	failed,
manteln	the mantle,mantle,
systematiska	systematic,systematical,
köra	run,drive,
koloniseringen	the colonization,colonization,
capitol	capitol,
dödsoffer	casualty,death victim,victim,
biskop	bishop,
krigsmakten	armed forces,
körs	driven,running,being driven,
birmingham	birmingham,
utrotning	extinction,extermination,
valutan	currency,
kommunal	communal,municipal,
döda	dead,
givit	gave,
matteus	matthew,matteus,
han	he,
grafit	graphite,
vetenskapsmän	scientist,scientists,
bnp	gdp,gnp,
fysikaliska	physical,
muhammeds	mohammed's,muhammad,muhammed's,
huvud	head,main,
hette	name was,named,
lunginflammation	pneumonia,
har	is,has,have,
hat	hatred,
hav	seas,sea,ocean,
präst	priest,
underliggande	underlying,
svensson	svensson,smith,
narkotika	drug,narcotics,
livsstil	life style,lifestyle,
dagar	says,day,days,
melodifestivalen	music festival,eurovision song contest,
uppmärksammade	observed,noted,noticed,
county	county,
bobby	bobby,
sedlar	bills,
alice	alice,
konsert	concert,
residensstad	city of residence,county seat,
sebastian	sebastian,
ola	ola,
old	old,
företräder	preferred trades,representing,
people	people,
reagera	reacting,reaching,
parlamentarisk	parliamentary,
delade	shared,divided,split,
kulmen	culmination,the acme,peak,
fot	foot,ft,
for	for,
varierande	variable,varied,varying,
fox	fox,
princip	principle,principal,
utser	chooses,appoints,
utses	is appointed,designated,appointed,
akademi	academy,
idéer	ideas,
myndigheter	authorities,agencies,
annan	another,
neptunus	neptunes,neptune,
stefan	stefan,
påminner	reminds,out,
hörde	heard,
binder	bind,tie,
olympiska	olympic,
möjligheterna	possibilities,the possibilities,
myndigheten	the authority,authority,
annat	alia,other,other; another,
evangelierna	gospels,the gospels,
army	army,
o	oh,
mynnar	opening,
klubben	club,
stjärna	star,
misstänkt	accused,suspect,suspected of,
nixon	nixon,
tillverkare	producer,manufacturer,
hänt	suspension,happened,
delvis	partial,partly,partially,
döpte	renamed,
psykiska	psychic,mental,
marshall	marshall,
som	as,which,
sol	sun,
lagliga	legal,lawful,
son	son,
psykiskt	psychic,mentally,
fci	fci,
delarna	the parts,parts,
artikeln	the article,
hantera	handle,
nova	nova,
säkerhetspolitik	safety policy,security,security policy,
joseph	joseph,
homo	homo,gay,
fria	free,
jane	jane,
 mm	millimeter,
happy	happy,
saltkråkan	salt crow,
jönköpings	jönköpings,
offer	victims,victim,
öppen	open,
förhållandet	the ratio,the relation,relationship,
förhållanden	relationships,conditions,n/a,
öppet	open,
verde	verde,
tigern	tiger,the tiger,
avsevärt	substantially,considerably,
förväntningar	expectations,
drabbat	affected,
gymnasiet	high school,gymnasium,
drabbar	affect,troubles,afflict,
polska	polish,
syften	purpose,
pest	plague,
syftet	purpose,
fansen	fans,the fan,
moderna	modern,
liberal	liberal,
föregångare	predecessor,precursor,
konung	king,
lunds	lund,lund's,
låtar	songs,
modernt	modern,
krävde	demanded,
ericsson	ericsson,
astronomiska	astronomical,
huvudperson	main person; main character,protagonist,main character,
dotter	daughter,
protester	protests,
läste	read,
republik	republic,
roll	role,
olja	oil,
reggae	reggae,
avskaffades	was abolished,abolished,
bostadsområden	residential,housing,residential areas,
palme	palme,
blått	blue,
vintrarna	the winters,winters,
modell	model,
rolling	rolling,
utbildade	educated,formed,
danske	danish,dane,
aragorn	aragorn,
tävling	competition,contest,
danska	danish,
sällan	seldom,rare,
povel	povel,
laddade	charged,
perioden	period,time,
kategorifödda	category born,category: born,
brasilianska	brasilian,brazilian,
trettio	thirty,
herren	lord,the lord,
perioder	periods; episodes,period,periods,
time	time,
erkända	acknowledged,recognized,
skatt	tax,
erkände	confession,acknowledged,
oss	center,us,
ost	cheese,
uppgifter	information,tasks,data,
stödjer	support,supports,
avalanche	avalanche,
uppgiften	the task,task,
atombomben	atomic bomb,the nuclear bomb,
stålgemenskapen	steel community,
inkomst	income,
behåller	retain,keeps,
machu	machu,
vet	know,
fängelset	prison,
intresserade	interested,
grön	green,
vem	who,
framställa	represent; depict; produce,produce,the installation,
bosnien	bosnian,bosnia,
musikstilar	music genres,music,
individer	individuals,subjects,
choice	choice,
individen	the individual,individual,
framställs	is depicted,prepared,
kombinerade	combined,
kusterna	the coasts,coasts,
initiativ	initiative,
lägre	lower,
inhemska	native,
energin	the energy,energy,
oppositionen	opposition,
team	team,
uppskattningsvis	estimated,approximately,an estimated,
årig	year old,minor,
jämnt	even,evenly,
nybildade	newly formed,newly established,
scen	scene,stage,
jämna	even,
fontsizes	fontsizes,
firandet	celebrate,the celebration,
måne	moon,
greve	count,earl,
känd	known,unknown,famous,
elton	elton,
köp	purchase,
kör	run,
kunskapen	the knowledge,knowledge,
beskydd	conservation,protection,
axel	axel,
bosatte	settled,
kön	gender,sex,
kunskaper	knowledge,
bosatta	residents,settled,
kusten	the coast,coast,
katter	cats,cat,
berättelsen	story,the story,
provinserna	provinces,the provinces,
galileo	galileo,
vintertid	winter-time,winter,
budskapet	the  message,the message,message,
katten	the cat,cat,
huvudsakliga	main,
studien	study,the study,
genomgående	consistently,through,pervading,
hälft	half,
bokstav	character,letter,
landslag	national team,
studiet	study,the study,
studier	studies,
love	love,
engelske	british,the english,english,
styrkan	strength; unit; force,strength,
publicera	publish,
kommit	to be,come,
presenterade	presented,
canis	canis,
sprids	spreading,spreads,
samlat	collected,single,gathered,
samlar	collect,salmar,collectors,
positiva	positive,
änglar	angels,
vuxna	adult,
sprida	spread,
judarna	the jews, therefore,jews,
positivt	positive,
samlag	intercourse,
effektiv	effective,
ställt	taken,put,set,
ställs	is,
dagars	day's,day,days,
relationerna	the relationships,relations,
tillträdde	assumed,took,
ställe	stalle,place,
hål	hole,hal,
ställa	make,set,installation,
tabellen	table,the chart,table; list,
dålig	poor,
grönt	green,
straffet	penalty,the punishment,
mörker	dark,darkness,
kunskap	knowledge,
gröna	green,
phoebe	phoebe,
påvisa	detection,show,prove,
stigande	rising,up,
locka	attract,tempt,
missförstånd	misunderstanding,misunderstandings,
locke	locke,
släktskap	relationship,kinship,
inkluderade	included,
rädda	save,lot of,
porträtt	portraits,portrait,
utnyttjade	utilized,used,
drama	drama,
milda	mild,
årligen	annually,yearly,annual,
skikt	layers,layer,
svenskan	swedish,the swede,
storleken	size,
trigonometriska	trigonometric,
européer	europeans,
levande	live,
riksdagen	parliament,the parliament,
gigantiska	gigantic,giant,
kungens	king,the king's,
löpande	running,assembly,conveyor (belt),
svart	black,
nyligen	recently,
data	data,
epost	e-mail,email,
portugisiska	portuguese,portugese,
stress	stress,
natural	natural,
bergarter	rock types,minerals,rocks,
undervisning	teaching,education,
påstod	claimed,said,
ss	ss,
sr	sr,
sv	sw,south west,
vikt	weight,
st	saint,
sk	so called,known,
so	so,
sm	s-m,swedish championship,
sa	said,
vika	fold,
se	see,
resulterar	resulting,result,results,
allvarliga	serious,severe,
resulterat	resulted,resulted in,
professorn	professor,the professor,
kong	(hong) kong,kong,
antingen	presumably,either,
allvarligt	serious,severe,
clinton	clinton,
irländsk	irish,ireland,
torg	square,
ingvar	ingvar,
dialekter	dialects,
utsätts	exposed,
torn	tower,
tilldelats	assigned,awarded,
turnera	tour,
museu	museum,
ersätts	replaced,
faderns	his father,the father's,
monopol	monopoly,
personlig	personal,
britter	britons,
hos	in; with,with,of,
änden	end,spirit,
öppnades	were opened,was opened,opened,
äldste	elders,eldest,
musiken	the music,music,
äldsta	oldest,
matcher	matches,games,
nation	nation,
records	records,
matchen	the game,match,
kategoripersoner	category of persons,
kantoner	cantons,
kravet	requirement,the demand,
twilight	twilight,
musiker	musicians,musicants,
atmosfär	atmosphere,atmospheric,
lockar	attracts,curls,
förväxlas	mixed up (with),confused,mistaken,
sidor	pages,sides,
säga	say,
skivkontrakt	record deal,record contract,
dominerar	dominate,dominates,
domineras	dominated,
runstenar	runestones,rune stones,
sägs	said (to be),said,
dominerat	dominated,
födelsedag	birthday,
prisma	prism,prisma,
dynamiska	dynamic,
greker	greek,greeks,
delstaterna	states,
förstöra	destroy,ruin; destroy,
väljas	elected,be elected,choose,
hinduer	hindu,hindus,
krav	requirement,conditions,demands,
kött	meat,cones,
riktigt	real,right,
ockupationen	the occupation,occupation,
specifikt	specifically,
sjuka	disease,sick,
densitet	density,
riktiga	real,
bränder	fires,
internet	internet,
roterar	rotates,
bla	blah,among others,
sfären	spheres,sphere,
garantera	ensure,guarantee,
vård	vard,nursing,healthcare,
våra	our,
singlar	singles,
sålde	sold,
bytt	changed,traded,switched,
byts	changed,replaced,
sålda	sold,salda,
väster	west,
vårt	our,each,
pilatus	pilatus,pilate,
dramaten	dramaten,
byte	change of,bytes,
byta	switch,change,trade,
föreställning	performance,
fyllt	filled,
pund	pound,
artister	artists,performers,
punk	punk rock,punk,para,
flandern	flanders,
solna	solna,
artisten	the artist,artist,
gordon	gordon,
startade	started,
givits	given,
jakob	jakob,
förmån	benefit,advantage; in favor of; benefit,
hård	diffcult,hard,
potter	pots,potter,
one	one,
slutet	end,
tsunamier	tsunamis,
hårt	hard,resin,difficult,
open	open,
ont	bad,
urin	urine,
city	city,
kraftigare	greater,more powerfully,
flytande	floating,liquid,
teologi	teology,theology,
skådespelarna	actors,
råolja	crude oil,
intill	beside,adjacent to,adjacent,
sjö	naval,lake,
nästa	next,
williams	williams,
animerade	animated,
vilka	who; which; that,who,which,
tillräckligt	sufficient,
irakiska	iraqi,irakish,
tillräckliga	insufficient,sufficient,
svenskarna	the swedes,swedes,
yttersta	furthest,supreme,highly,
provins	province,
dygn	day,
fiskar	fishes,fish,
uppenbarelser	revelations,
berlinmuren	berlin wall,the berlin wall,
kamprad	kamprad,
motståndarna	the opponents,opponents,
tankar	tank,thoughts,
sak	thing,matter; case,substance,
san	san,
sam	co,
generation	generation,
konsekvenser	consequences,
argument	arguments,argument,
församlingar	parishs,assemblies,
say	say,
känslan	feeling,the feeling,sense,
burundi	burundi,
allen	allen,
utgåva	edition,issue,
staden	city,the city,
priserna	prices,the prices,
skickades	was sent,sent,
takt	rate,
general	general,
styrelsen	the board,board,
zoo	zoo,
jefferson	jefferson,
massa	mass,
övrigt	other,
förändringen	the change,change,
föder	give birth,gives birth,give birth of,
muslimer	muslims,
finlands	finland's,finlands,
sekreterare	secretary,
tränare	coach,
mynt	coins,coin,
religionen	religion,the religion,
betyda	mean,
religioner	religions,
forskningen	the science,research,
rådets	council,
kontroversiell	controversial,
driva	operate,run,
förändras	changes,
inledningen	introduction,the beginning,the introduction,
ursprung	origin,root,
fredspriset	nobel peace prize,peace price,peace prize,
rykte	reputation,
färdig	pre,done,
katekes	catechism,
rött	cane,red,
olagligt	illegal,
axl	axl,
genomförts	out,
beckham	beckham,
vart	each,
ledd	led,
dimensioner	dimensions,
dahléns	dahlens,dahlén's,dahlen,
sjöss	sea,
antalet	number,the number,
stärkte	strengthened,increased,
slog	hit,
hockey	ice hockey,hockey,
caroline	caroline,
carolina	carolina,
belgien	belgium,
kategorimusik	category music,
återvänder	returns,atervander,
inlägg	post,
beatrice	beatrice,
egentliga	real one,actual,
platta	flat,
undersöka	study,understand,research,
rörande	concerning,
spetshundar	tip of dogs,
ländernas	countries',the countries,countries,
artist	artist,
råd	advice,council,
enighet	unity,
översättningen	translation,the translation,
roger	roger,
ljudet	the sound,noise,
varna	varna,alerting,
sträcka	distance,
monark	monarch,
erbjöds	offered,
dagsläget	present situation,current situation,
hämtar	download,is,gets,
spetsen	edge; top,tip,
brännvin	schnaps,aquavit,
snabbare	rapid,faster,
behovet	need,the need,
up	i[,up,
nederbörden	precipitation,the precipitation,
skärgård	archipelago,cutting garden,archipelagos,
talman	spokesperson,president,speaker,
ordspråk	saying,proverb,proverbs,
enhetlig	single,unitary,uniform,
utgörs	consists of,is,make up,
förvaltning	management,administration,
källa	source,
kritiserade	critisized,criticized,criticised,
begränsningar	limitations,limits,
upplever	experiencing,experience,
kontrakt	agreement,contract,
utgöra	compose,make up,
kilometer	kilometer,kilometers,
revolutionär	revolutionary,revolutions,
små	small,little, small,
gäller	of,refer to,grating,
amerikanskt	american,
anledningarna	reasons,the reasons,
söka	search,searching,
screen	screen,
fynd	finding; finds,findings,
antika	ancient,
amerikanske	american,the american,
awards	awards,
inverkan	impact,influence,effect,
amerikanska	u.s.,american,
mariette	mariette,
basisten	bassist,basist,the basist,
skönlitteratur	nonfiction,fiction,
mans	man's,
nationell	national,
erics	erics,
rekord	record,
mani	mani,mania,
tillsätts	added,appointed,appoints,
långsammare	more slowly,slower,
upproret	the upprising,revolt,rebellion,
klimat	climate,
hamnade	landed,ended up,
anta	assume,assume; adopt,adopting,
drogs	was pulled,was,
därtill	thereto,
teddy	teddy,
farfar	paternal grandfather,grandfather,
west	west,
airlines	airlines,
bolag	company,
luft	air,
cupen	the cup,cup,
lidit	sustained,suffered,
lånat	borrowed,
förr	sooner; past,sooner,before,
formen	the form,form,
formel	formula,
sångerska	songstress,singer,
regimer	regimens,regimes,
warhol	warhol,
tillåter	allows,allow,
tillåtet	allowed,
pernilla	pernilla,
former	forms,
landskapen	the landscapes,landscapes,landscape,
samling	concentration,collection,
representativ	representative,
landskapet	landscape,
värderingar	evaluations,values,
situation	situation,position,
föregångaren	predecessor,it's predecessor,
peruanska	peruvian,peruan,
aborter	abortions,
aluminium	aluminum,
startar	begins,start,starts,
bror	brother,
ekonomi	economic,economy,
tillåtelse	permission,allowed,
sammanfaller	coinciding,coincides,
beteckna	denote,
ohälsa	disorders,
världsbanken	world bank,
undersökning	study,survey,
träffat	met,
ärftliga	genetic,
otto	otto,
träffas	reached,meet,
oceanen	the ocean,ocean,
ekologi	ecology,
ludwig	lugwig,ludwig,
nationalparker	national parks,
singapore	singapore,
sägas	is said,is said (to be),said,
lindgrens	lindgren's,lindgrens,lindgren,
följer	resulting,
förkortning	abbreviation,
senator	senator,
dsmiv	dsm-iv,
personlighetsstörning	personality disorder,
måla	target,
tillfälle	instance,time,occasion,
gestalter	beings,figures,
avser	regards,regard,refers to,
avses	refered,regard,referred,
ifrågasatt	question,questioned,
iraks	iraq,
gudomliga	divine,
summer	sommar,
förluster	loss,losses,
bokförlaget	bokförlaget,publisher,publishing house,
berättelse	tale,story,'s re,
rest	remain,residual,rest,
koncentration	concentration,
spårvagnar	trams,
psykologisk	psychological,
likheter	similarities,similarity,
resa	travel,
libyen	libya,
förlusten	loss; defeat,loss,
avbryta	cancel,
judarnas	jews,
kastar	throws,to throw,
heliga	saints,holy,holy; holy,
unika	unique,
sprider	spreads out,spread,spreads,
helige	holy,
miljon	one million,million,
instrument	intrument,
fördrevs	was banished,ford described,driven away,
sänka	lower,
infördes	introduced,
unikt	unique,
heligt	holy,heligit,
störst	most,
snart	soon,once,
vinkel	angle,
dark	dark,
regim	regimen,regime,
unesco	unesco,
litteraturen	literature,
skadade	wounded,damaged,
stammar	strains,stutters,tribes,
statsreligion	state religion,
framsteg	progress,
tvserie	tv serial,
carl	carl,
tsunami	tsunami,
ekonomier	economies,
stupade	fallen,killed,
fossila	fossilized,fossil,
inter	inter,
intet	nothing,no,
jobbar	work,does the work,
nämnas	mentioned,worth mentioning,include,
what	what,
domkyrkan	cathedral,the cathedral,
ursprungsbefolkning	native population,indigenous,
ekman	ekman,
kännedom	known,knowledge,
närheten	near,the vicinity,
björn	björn,bear,
föreslog	suggested,propose,
institutionerna	institutions,
ddr	ddr,
än	than,yet,
exil	exile,
inkluderar	include,includes,
cannabis	cannabis,
varsin	(one) each,opposite,
är	is,
atomkärnor	nuclei,nuclear particles,atomic cores,
ingående	input,enter into,in depth,
västerås	vasteras,västerås,
katolsk	catholic,
långstrump	longstocking,
jacksons	jackson's,jacksons,jackson,
nivån	level,
medlemsstater	member,member states,member-state,
stone	least,
organisationen	organization,the organization,
ace	ace,
herrlandslag	men's national team,women's national teams,
vissa	some,
populationen	the population,population,
befinner	is,placed; situated; positioned; are,
digerdöden	black death,the black death,
populationer	populations,
lyssnade	listened,
organisationer	organizations,organisations,
industri	industry,industrial,
visst	specific,certain,
regissör	director,
berger	berger,
upplevelser	experiences,
ronden	round,
bryts	breaks,
nationalencyklopedin	national encyclopedia,the national encyclopedia,
image	image,
säkerhetsrådet	security,
partiet	the party,portion,
bryta	break,
partier	portions,parties,
angola	angola,
bergen	the mountains,mountain,mountains,
het	hot,up to date,
företag	company,companies,business,
kallats	was called,called,
förintelsen	holocaust,the genocide,
philadelphia	philadelphia,
evangeliska	evangelical,
söker	searches,seek,seeks out,
hel	full,(whole) lot (of),
hem	home,back,
hamnen	harbour,the harbour,
sover	sleep,
enorm	huge,enormous,
hänger	depends,hanger,
hänvisning	reference,
project	project,
dagen	day,
complete	complete,
hells	hells,
bevarat	preserve,preserved,
bevaras	are protected,preserved,
mick	microphone,mick,mike (microphone),
kontroverser	controversies,contraversies,
språkliga	linguistic,
bevarad	kept,preserved,
åttonde	eighth,the eighth,
rush	rush,
sällskap	company,groups,
jamaicas	jamaicas,jamaica's,
hexadecimalt	hexa-decimal,hex,
kvartsfinalen	quarter finals,quarterfinals,
utmed	along,
vinkeln	angle,the angle,
afrodite	aphrodite,afrodite,
förbundsstat	federal,federal state,
produkt	product,
puls	pulse,
krona	crown,
ac	ac,
ab	ab,
brodern	the brother,brother,
johnny	johny,johnny,
redovisas	reported,shown,accounted for,
gustafs	gustafs,gustaf's,
am	am,
al	alder,
bronsåldern	bronze age,the bronze age,
as	as,
beordrade	commanded,ordered,
övernaturliga	supernatural,over natural,
av	of,
håll	ways,hold,
väsentligt	substantially,relevant,
testamentet	testament,
vore	would,were,
federala	federal,
rökning	smoking,
utförde	did,
svårt	hard,difficult,
belönades	rewarded,awarded,
isolerad	isolation,isolated,
svåra	answering,difficult,
avslöjade	revealed,
såsom	such as,like,
gifta	marry,married,
värt	worth,
koppar	copper,
gifte	married,
medverkan	the contribution,participation,
kvarstod	remained,
kategorisvenskspråkiga	category swedish-speaking,
terra	terra,
medverkat	participated,
medverkar	contributes,contribute,
terry	terry,
vanliga	ordinary,regular,usual,
forntida	pristine,ancient,prehistoric,
kommunen	municipality,
skador	damage,
århundradena	centuries,
beteckning	indication,label,
adam	adam,
omgivningen	surroundings,the surrounding,ambient,
decennierna	decades,the decades,
original	original,orignal,
renässans	renaissance,
känslor	music,feelings,
släppt	self-indulgent,relinquished,released,
släpps	released,(is) released,
elektron	electron,
halsen	throat,the neck,the throat,
anpassning	adaption,adjustment,
myntade	coined,
års	years (age),year,years,
släppa	release,
likartade	similiar,similar,
 kmh	km/h,
norr	north,
skogarna	the forests,forests,
number	number,
pojkvän	n/a,boyfriend,
ullevi	ullevi,
tv	tv,
romanen	novel,
nederbörd	rainfall,precipitation,
to	to,
mildare	cooler,milder,mild,
romaner	novels,
th	th,
nord	north,
te	tea,
sättas	turn,added,
ta	to,take,
avlägsna	distant,remove,
använder	using,uses,
arvet	the inheritance,heritage,
telefonen	phone,the telephone,
strand	beach,
utländsk	foregin,foreign,
sant	true,
ensamma	alone,
djurarter	species of animals,animal species,species,
borrelia	borrelia,borreliosis,
muslimska	muslim,
utsåg	declared,appointed,
sand	sand,sandy,
siffrorna	figures,the numbers,numbers,
områdets	the area's,of the area,area,
harry	harry,
sann	true,
språkbruk	language (use); parlance; phraseology,parlance,language,
förmedla	pass; express; mediate,pass,
döttrar	daughters,
samoa	samoa,
påståenden	claims,assertions,
synd	sin,
dödsstraff	death penalty,
utökade	expanded,increased,
vägnät	network,
pass	an,
givaren	donor,the giver,dealer,
syns	seen,visible,
richard	richard,
stängt	closed,
delen	part,
soldater	soldiers,
islams	islams,islam's,
leif	leif,
gjorts	made,done,
hänsyn	light,consideration,
full	full,
gruppen	the group,group,
själen	soul,the soul,
arkeologiska	archaeological,
november	november,
legend	legend,
motstånd	resistance,opposition,
äventyr	adventure,adventures,
hindra	hinder,prevent,stop,
traditionella	traditional,conventional,
exklusiv	exclusive,
traditionellt	traditional,
social	social,
action	action,
oftare	more often,more frequently,more,
varelser	creatures,
medlemskap	membership,
kommunistpartiet	communist party,the communist party,
vid	in,by,at,
ordinarie	permanent,ordinary,regular,
vii	vii,
vin	whine,wine,
young	small,
juridiskt	legally,juridical,judicial,
vis	vis,wise,way,
kuiperbältet	the kuiper belt,the cuyper belt,
vit	white,
spelaren	the player,
motsatsen	the opposite,opposite,
biskopen	bishop,the bishop,
mors	mother,mothers,
petroleum	oil,petroleum,
underordnade	subordinate,subordinates,
pearl	pearl,
sitter	is,serve,sit,
presenterades	presented,
rhen	the rhine,rhine,
dödligt	lethal,deadly,
mora	mora,
bevis	certificate,evidence,
mord	murder,
ragnar	ragnar,
uppskattad	estimated,appreciated,
berättade	told,
uppskattas	is appreciated,estimated,appreciated,
uppskattar	estimated,estimates,
schweiz	switzerland,
undergång	during navigation,doom,destruction,
socialt	socially,social,
inträffade	occurred,happened,
medelklassen	middle class,
science	science,
monoteistiska	monotheistic,
klp	klp,
sociala	social,
morgan	morgan,
kapitalism	capitalism,
studenter	students,
läkaren	the doctor,physician,
samväldet	commonwealth,the commonwealth,
nobelpriset	the nobel prize,nobel award,
säljas	is sold,sold,
nordvästra	northwest,north western,
skadliga	harmful,deleterious,
huvudstaden	capital,
mellersta	middle,the middle,
states	states,
stater	states,
spansk	spanish,
järnvägsnätet	railroad network,rail,
information	information,
vägnätet	road network,
uteslutande	exclusivly,only,exclusively,
hugo	hugo,
uppfattade	perceived,perceive,
ansetts	considered,regarded,regarded; viewed (as),
uppnått	met,achieved,
lejon	lion,
riksdagens	the parliament's,the parliaments,
retorik	rhetoric,
variant	variant,type,variety,
hustru	wife,
produktionen	production,the production,
referens	reference,
lanka	lanka,(sri) lanka,
köpte	purchased,bought,
barnens	the child's,childrens,
komplext	complex,
anklagade	accused,
pucken	the puck,
komplexa	complex,
utvidgning	enlargement; expansion,enlargement,
hållit	held,maintained,kept,
nationerna	the nations,nations,
blommor	flowers,
trade	esterified,
östblocket	east block,the eastern bloc,cheese block,
scott	scott,
kvinnors	women's,women,
aktiviteter	activities,activity,
anställda	employed,
radion	the radio,radio,
vietnamkriget	the vietnam war,vietnam war,
känsla	feeling,sense,
alla	all,everyone,
högskola	college,
protestanter	protestants,
caesars	caesars,
miljön	environment,the environment,
termen	the term,term,
filip	phillipe,filip,
termer	term,terms,
allt	all,
alls	all,
få	have; make; few,gain,fa,
van	van,
isaac	isaac,issac,
konstruerade	constructed,
samhällets	society,of society,
berömda	famous,
inleda	initiate,
källan	source,kallan,the source,
beräkna	calculated,calculate,
privilegier	privileges,
inledande	initial,
produceras	produced,
producerar	producing,produces,
grekisk	greek,
producerat	produced,
introducerade	introduced,
producerade	produced,
olycka	incident,accident,disaster,
intåg	entry,advent,
budskap	message,
målning	painting,
graviditet	pregnancy,
blodet	the blood,blood,
denne	his,that he,he,
denna	that,
härrör	derived,
enstaka	occasional,single,
england	england,
populärt	popular,popularly,
sydöst	south east,southeast,
doser	dose,
populära	popular,
blues	blues,
förespråkade	advocate,advocated,
kretsen	the order,circuit,
finner	found,finds,
uppfördes	was constructed,built,constructed,
återkomst	return,
omröstningen	vote,the election,
kopplad	connected to,connected,
garvey	garvey,
avgick	resigned,retired,
research	research,
norska	norwegian,
uppstått	resulting,arised,arisen,
sammanfattning	summary,
besökte	visited,
kopplat	coupled; connected,connected,coupled,
hallucinationer	hallucinations,
highway	highway,
medel	middle,medium,
sparken	park,gets fired,fired,
alltmer	increasingly,more and more,
stjärnor	stars,
poeter	poets,
driver	driver,run,drive,
båda	both,
både	both,
kostade	cost,
ålands	Åland island's,the Åland island's,aland,
kärnkraft	nuclear power,nuclear,
poeten	poet,the poet,
teknologi	technology,
definition	defined,definition,
service	service,
turistmål	tourist destination,tourist attraction,
hjärta	heart,
naturens	nature's,nature,
samlas	together,
omfattar	encompass,include,
skolan	school,
w	w,
nivåer	levels,
besök	visit,
uppenbarelse	apparition,revelation,
principen	the principal,principle,
bidragit	contributed,
kristna	christian,
foten	foot,
skiftande	shifting,
spekulationer	speculation,speculations,
såg	see,saw,
gemensamma	joint,common,
avel	breeding,breed,
liknas	compared to,likened,
liknar	similar,similar to those,
tove	tove,
saint	saint,
sår	sir,wound,
missade	failed,
besläktat	related to,related,
läggas	laid,added,
chefen	head,commendant; commander,
tappade	lost,
zeus	zeus,
borgmästare	mayor,
moder	parent,mother,
svår	severe,difficult,
bidrog	contribute,contributed,
obama	obama,
organiseras	organizes,organized,
återkom	return,returned,feedback,
organiserat	structured,
niklas	niklas,
koncentrerade	concentrated,
marknadsekonomi	market,market economy,
freud	freud,
organiserad	organised,organized,
nikolaj	nikolaj,nicholas,
ägg	eggs,egg,
äga	be,own,aga,
väljer	select,elects,
inkluderas	include,is included,
statyn	the statue,statue,
generationen	generation,the generation,
förstörelse	destruction,
inkluderat	included,including,
ägt	taken,
generationer	generation,generations,
astronomin	the astronomy,astronomy,
visats	shown,demonstrated,
framåt	forward,forth,
varianten	version,variant,
norstedts	norstedt's,norstedts,collins,
kongokinshasa	kong kinshasa,democratic republic of the congo,congo kinshasa,
varianter	variants,varieties,diversities,
vinterspelen	winter games,
arabisk	arabic,
edison	edison,
sydostasien	south east asia,southeast asia,
brooklyn	brooklyn,
kväve	nitrogen,
plan	flat,level,
kombinationer	combinations,
arter	species,
utsattes	subjected,were exposed,exposed,
cover	cover,
kanalen	the channel,channel,
kanaler	channels,
monarki	monarchy,
arten	species,
kombinationen	the combination,combination,
golf	golf,
gold	gold,
omfattade	included,covered,
falska	false,
presidentens	the president's,president,the presidents,
detalj	detail,
karaktär	character,
falskt	false,
richmond	richmond,
framgångar	successes,success,
existensen	existence,
betydelser	values,meanings,
jämföra	compare,
befolkningstätheten	population density,n/a,state of the population,
wayne	wayne,
betydelsen	the meaning,significance,
jämfört	compared to last,compared,compared (to),
kontor	office,
karakteristiska	characteristic,
genomgick	underwent,
gratis	free,
evolutionen	evolution,the evolution,
tekniken	techinque,art,the technology,
tekniker	technician,
actress	actress,online,
utbildningen	education,
föll	fell,
erkännande	recognition,
victoriasjön	victoria lake,lake victoria,
tanken	the thought,idea,
ledare	conductors,leader,
cry	cry,
populärmusik	popular music,pop music,
byten	byte,
allmän	general,
river	tear,river,
sköt	shot,
någon	someone,anybody,
nietzsches	nietzsche,nietzsche's,
ses	be,are seen,
ser	see,sees,
koranen	the koran,the quran,
sex	six,
sed	sed,thirst,
psykologiska	psychological,
uppkomsten	onset,origin,
moçambique	mozambique,
järnväg	railroad,rail,railway,
sen	then,since,
något	any,something,
sorters	kinds of,kinds,
institutet	institute,the institution,
församlingen	parish,congregation,
påverkat	influenced,affected,
guinea	guinea,
neutralitet	neutrality,neutral,
fission	fission,
kejsarens	emperor,the emperor's,emperors,
stärkelse	starch,
alqaida	al-qaida,al-qaeda,
rita	paint,draw,drawing,
europe	europe,
europa	europe,european,
påverkar	affecting,
giftermål	marrige,marriage,
medveten	conscious,aware,
avvikelser	abnormalities,deviations,derivations,
medvetet	consciously,conscious,
fame	fame,
stadsdel	city district,neighborhood,district,
demografiska	demographic,demographical,
forskare	researcher,researchers,scientists,
bästa	the best,best,
medicinering	medication,
förändring	change,
bäste	best,
messias	messiah,
stå	stand,
halmstads	straw city,halmstad's,
kopia	copy,
samma	the same,same,
transeuropeiska	trans-european,transeuropean,
upprättades	was established,establish,
krisen	crisis,the crisis,
kriser	crises,
church	church,
allierade	allied,allies,
decennium	decade,
sommaren	summer,the summer,
pressfrihetsindex	press freedom index,pressfrihetsindex,
väntade	expected,expected; were waiting,waited,
tillväxt	growth,
potentiellt	potential,
kyrilliska	cyrillic,
upprättas	established,establish,
blod	blood,
pågår	(in) progress,underway,
föranledde	brought about,led,
beskrevs	was described,described,
skönhet	beauty,
östafrika	east africa,
fire	fire,
mind	mind,
fira	celebrate,
hovrätten	court of appeals,the court of appeal,
fritz	fritz,
uppleva	experience,
fritt	free,
föreningar	associations,organizations,compounds,
systematik	systematics,systematic,
handling	action,act,
framträder	stand out,stand,appear,
projekt	project,
budget	budget,
guldbollen	the ball,golden ball,guldbollen,
individerna	subjects,the individuals,
bestående	comprising,lasting,
brottslighet	criminality,crime,
pressen	press,the pres,
real	real,
föreställa	pretend; imagine,imagine,
arbete	work,work; labor,
vol	v,
von	von,
owen	owen,
motors	engine's,motor,
teoretisk	theoretical,
erkänna	recognize,
slöts	concluded,signed,
lokaler	facilities,studios,place,
korruptionsindex	corruption perceptions index,corruption index,
hovet	court,the court,
kritiker	critics,critiques,
barney	barney,
gärning	deed,
möjlighet	an opportunity,oppertunity,possibility,
omvandlas	convert,converted,
omvandlar	converts,transmuted,
skalet	shell,the shell,
tillkom	hold back,resided,
barnen	children,
arméer	armies,army,
kritiken	criticism,the criticism,the critique,
laddning	charge,
kategoriavlidna	category deceased,
snarare	rather,
republiken	the republic of,the republic,
republiker	republics,
skapade	made,created,
debatten	debate,the debate,
kring	on,around,
djurgården	djurgården,zoo,
fyra	four,
vargar	wolves,
euro	euro,
normala	normal,
krigsmakt	military power,armed forces,
person	person,
kelly	kelly,
johan	johan,
kontakter	contact,contacts,
finansiellt	financial,
nacka	nacka,
tunnelbana	subway,
stränder	beaches,
släppas	released,be released,
telegram	telegram,
stockholms	stockholm's,stockholm,
finansiella	financial,
kontakten	connector,conntact,the contact,
mandat	mandate,
fascistiska	fascist,fascistic,
rebecca	rebecca,
festivalen	festival,the festival,
symbolisk	nominal,symbolic,
nordväst	north west,northwest,
festivaler	festivals,
jönssonligan	jönssonligan,jonssonligan,
tomas	tomas,
hennes	her,
format	shaped,format,
turnéer	tours,
teologiska	theological,
melker	melker,
avvisar	reject,
skara	city in south-central sweden (uppland),crowd,
samarbete	collaboration,co,
ivar	ivar,
västsahara	western sahara,
samarbeta	collaborate,co,cooperate,
da	da,
talrika	numerous,
funnit	found,
skarp	sharp,crisp,
utlösa	trigger,
informationen	the information,
patrick	patrick,
ivan	ivan,
alexandra	alexandra,
ulrich	ulrich,
vojvodina	voyvodina,vojvodina,
lenin	lenin,
saknar	lacks,lack(-s),missing,
saknas	missing,
användbar	useful,
utvecklades	developed,(was) developed,
avskaffade	abolished,absolished,
nåd	mercy,grace,
wallenstein	wallenstein,
öka	oka,increase,increasing,
förtjust	fond,delighted,
trafiken	traffic,the traffic,
turnerade	toured,
religion	religion,
vacker	beautiful,
riksförbundet	national association,
säger	said,says,claims; says,
be	be,
norra	north,northern,
ugandas	of uganda,uganda,
västra	west,vastra,western,
bl	bl,short of "bland" - in the context: bl. a (bland annat) = among others,
vagnar	carts,wagons,carriges,
bo	living,
bk	bk,
plocka	pick,
engelska	england,english,
tid	time,
ordning	system,
santa	santa,
by	by,village,
källor	source,
ideologin	ideology,the ideology,
bosättningar	settlements,bosattningar,
soldaterna	soldiers,the soldiers,
dagligen	day,daily,
gemenskaperna	communities,community,
aggressiv	aggressive,
arméerna	armeerna,armies,
stuart	stuart,
fungerande	functioning,effective,working,
för	of,to; for,for,
papper	paper,
texterna	text,
inte	not,
inta	taken,
colorado	colorado,
syret	the oxygen,oxygen,
hemingway	hemingway,
efterföljande	subsequent,
spridas	spread,disseminated,
kraven	the demands,requirements,
popsångare	popsinger,pop singer,
uppkallad	named,
orsaken	reason,cause,
förlaget	publisher,the publisher,the publishing company,
seger	victory,
veckor	weeks,
kategorimusikgrupper	category of music groups,
dröja	take,
utbröt	erupted,broke out,
u+	u +,
samerna	sami,the lapp,
knuten	tied to,bound,knot,
hälften	the one half,half,
fattigdom	poverty,
förbindelse	connections,connection,
européerna	europeans,
poster	positions,post offices,
rörlighet	mobility,movement,
pastor	pastor,
begreppen	the concepts,the terms,terms,
begreppet	the term,term,concept,
posten	post,the position,
atom	atomic,atom,
kritisk	critical,
line	line,
lovade	promised,
lina	line,lina,
dröm	dream,syndrome,
fader	father,
cia	cia,
ut	out; up,out,
dom	judgement,conviction,
drogmissbruk	drug abuse, substance abuse, drug addiction,drug,
eddie	eddie,
us	oss,
ur	from,out,
konventionella	conventional,
distrikt	district,
uk	uk,
protestantiska	protestant,protestantic,
galaxer	galaxies,
testamente	testament,will,wills,
professor	professor,
översvämningar	flooding,floodings,
nämner	mentions,names,
spontant	spontaneous,spontaneously,
diverse	some,miscellaneous,
utbyggt	develpoed,built,extended,
makedonska	macedonian,makedonish,
nationalism	nationalism,
inblandning	involvement,incorporation,
matematiken	mathematics,
händelsehorisonten	event horizon,the event horizon,place else horizon,
räkna	count,special,
värld	world,
edwards	edwards,edward's,
são	sao,
skrivits	down,been written,
innehåller	include,contains,
nordafrika	north africa,
innehållet	content,contents,
matematiker	mathematician,
siffror	figures,numbers,
upplaga	edition,submission,
individuella	individual,
besegra	defeat,
dominerades	was dominated,dominated,
radikala	radical,
djurgårdens	djurgården's,
lucia	lucia,
ägnar	spend time,dedicated,spends time,
konstantinopel	constantinople,
riskerar	could,risks,there is a risk,
springsteen	springsteen,
radikalt	radical,radically,
slås	beat,is hit,slas,
alltså	so,therefore,really,
land	country,
passagerarna	passengers,the passengers,
uppträdande	performance,appearance,conduct,
symtom	symptoms,symptom,
age	do,age,
härstammar	derived,stems,
texten	text,the text,
sawyer	sawyer,
texter	texts,
majs	corn,
förväntas	expected,
persbrandt	persbrandt,
släpptes	released,was released,
alltför	all too,way too,exessive,
bakåt	backwards,reverse,
anorektiker	anorectics,anorexic,anorectic,
turkisk	turkish,
dyraste	most expensive,
hamnar	lands,ports,
hamnat	got,ended up,got in to,
listade	listed,
dickinson	dickinson,
dancehall	dance hall,dancehall,
sent	late,
garden	garden,
märken	brands,sign,
kedjan	chain,the chain,
palestinier	palestinians,palestinian,
kommunistiska	communistic,communist,
flöde	feed,
drogen	the drug,drug,
vinner	gaining,wins,win,
känner	knows,know,
överleva	survive,survival,
tillhörande	associated,belonging to,belonging (to),
magic	magic,
tro	believing,think,
påverka	impact,influence,
harbor	harbor,
eva	eva,
tre	three,
jobbet	work,the job,
romerska	roman,
överlevt	survived,
romerske	roman,
opinionen	opinion,
agera	act,
leonardo	leonardo,
bolsjevikerna	bolsheviks,the bolsheviks,
natur	nature,
regelbundna	regular,
ställde	set,stood up,asked,
årtionden	decades,
video	video,
förhållandevis	relatively,
förkortningar	abbreviations,
legitimitet	legitimacy,
victor	victor,
antog	adopted,
index	index,
expressen	expressen,
anton	anton,
praktiken	effectively,practice,practically,
indiens	india's,indias,
suveräna	terrific,supreme,sovereign,
möjliggör	enables,enable,
birk	brik,birk,
indian	indian,
ledande	conductive,leading,
wembley	wembley,
stadskärna	city core, city center,town,town centre,
led	suffered,step,
lee	lee,
lyckades	managed,succeeded,
upphovsrätten	copyright,
sålunda	thus,
leo	leo,
les	les,
let	cleanly,
lev	live,lev,
hälsa	health,tell (him i said hi),
talang	talent,
begravd	buried,
motorvägarna	highways,the highways,
tegel	brick,
casino	casino,
titanic	titanic,
förutsätter	assume,requires,assumes,
högste	supreme,highest,chief,
insulin	insulin,
högsta	highest,
opinion	opinion,
sekel	centuries,century,
huvudvärk	headache,
emot	vis,against,
förlora	lose,
oxenstierna	the oxenstierna,oxenstierna,
mening	meaning,meanings,sentence,
fotosyntesen	photosynthesis,
anatolien	anatolia,
andreas	andreas,
varmare	heater,warmer,
sekulär	secular,
illegal	illicit,illegal,
hemlig	secret,
elever	students,
godkänna	approve,
klaviatur	keyboard,
toy	toy,
orkester	orchestra,
projektet	project,
herbert	herbert,
existerade	existed,existing,
författning	constitution,
samspel	interaction,teamwork,
ytterst	very; extremely,highly,
överlevande	survivors,survivor; survivors; surviving,
villor	houses,villas,
edwall	edwall,
lokalt	locally,local,
nordliga	northernly,northern,
advokat	bar,lawyer,
ortodoxa	orthodox,
lokala	local,
peka	point (at; to; in),point,
gustafsson	gustafsson,
upprätthålla	maintain,keep up,maintaining,
process	process,
artiklar	items,
etta	number one,first,one,
tryckta	printed,
high	high,
syre	oxygen,
hercegovina	herzegovina,
sydöstra	the southeast,south east,south eastern,
föregående	preceeding; previous,previous,
halmstad	halmstad,halmstad's,
gitarr	guitar,guitarr,
saknade	lacked,missed,missing,
delad	shared,divided,
västerbottens	västerbottens,västerbotten's,west bothnia,
latinska	latin,
hormoner	hormons,hormones,
delas	shared,divided,
delar	proportions,parts,
delat	shared,divided,
sydvästra	southwest,southwestern,
kriminella	criminal,
gunwer	gunwer,
amerika	american,america,
djurens	the animals,animal,
profeten	prophet,the prophet,
insatser	action,
regeringsmakten	govermental power,government power,
platt	flat,plate,
democracy	democracy,
väckt	brought,awaken,woken,
slutsatser	conclusions,
frågor	questions,
element	elements,
lundgren	lundgren,
nancy	nancy,
napoleons	napoleon,napoleon's,
byggnadsverk	building,construction,edifice,
borde	should,
handboll	handball,
diskar	disks,
houston	houston,
möjligt	possible,
hårdast	the most,the hardest,hardest,
universiteten	universities,the universities,
frånvaro	absent,absence,
hunnit	reached,had,had time to,
universitetet	the university,university,
bensin	gasoline,
sydligaste	southernmost,most southern,
möjliga	possible,
solvinden	the solar wind,solar wind,
övergrepp	assault,abuse,assult (-s),
eliten	the elite,elite,
uppdelat	divided,split,
fristående	independent,stand-alone,
tecknet	the sign,sign,
uppdelad	divided,split,
puerto	puerto,port,
beståndsdelar	constituents,elements,
ovanlig	unusual,rare,uncommon,
konkurs	bankrupcy,bankruptcy,
bekant	known,acquaintance,
bryter	breaks,breaking; violating,
hemmaplan	home,home turf; domestic (level),
dock	nevertheless,however,
utgår	deleted,
rotation	rotation,
huvuddelen	bulk,main part,
sönder	broken,probes,
orange	orange,
peking	beijing,peking,
välfärd	wealth,welfare,
intressen	interests,
fortsätta	remain,continue,
smallwood	small wood,smallwood,
burton	burton,
books	books,
intresset	interests,the interest,interest,
frac	fraction,
bay	bay,
etymologi	etymology,
matrix	matrix,
borderline	borderline,
billiga	cheap,
utbildad	educated,formed,
enskilda	individual,
anledningen	reason,therefore,
umgänge	company,intercourse,
kapitalismens	capitalism's,capitalism,
marxistiska	marxist,
bekräftades	confirmed,was confirmed,
fram	until,out,
undertecknades	signed,
legat	formed,layed,
redskap	device,tool,
egenskaperna	the qualities,properties,
mötte	motte,met,
kalle	kalle,
påverkats	influenced,affected,
melankoli	melancholy,
uppe	top,up,(on) top, up, above,
lundin	lundin,
förts	brought,cont,
tempererat	temperate,tempered,
dubbel	double,
liggande	placed,overhead,lie,
kompositör	composer,
krävt	taken,required,
våldsam	violent,
krävs	needs,required,requires,
david	david,
blanda	mix,
profeter	prophets,profets,
krets	sphere,circuit,
helst	rather,anyone,any time,
davis	davis,
hussein	hussein,
kräva	require,demand,
skillnad	difference,unlike,
playstation	playstation,
åring	year old,years,
komplicerade	complex,
jesus	jesus,
användningsområden	possible use,applications,
schweiziska	swiss,
muhammad	muhammad,
nordkoreanska	north korean,
studerade	studied,
nationalistiska	nationalist,nationalistic,
festival	festival,
system	system,
bygget	the construction,construction,
syster	sister,
hebreiska	hebrew,
tränga	push (aside),cut in,permeate,
teatern	the theater,theater,
blivit	become,was,
utbyggnad	development,addition,expansion,
havet	sea,
pristagare	laureate,prizewinner,
konservativ	conservative,
utländska	foreign,
haven	the seas,
visdom	wisdom,
hampa	hemp,
samverkar	co,co-operating,co-operates,
roberto	roberto,
stewie	stewie,
roberts	roberts,
reagans	reagan's,reagan,
troende	believers,faithful,
vecka	week,
jonatan	jonatan,jonathan,
räcker	enough,sufficient,
användaren	the user,user,
inre	inner,
förslag	proposal,'proposal,proposed,
flygplats	airport,
kritiskt	critical,
instruktioner	instructions,
mills	mills,
filosofin	philosophy,the philosophy,
sinatra	sinatra,
sekvens	sequence,
kritiska	critical,
best	best,
uppträdde	appeared,perform,occurred,
viss	certain,some,
finsk	finnish,
slutsatsen	concluded,the conclusion,
säkert	securely,
när	when,
nät	web,net(work),
minoritet	minority,
detta	this,that,
vardagen	the weekday,everyday life,
kvinnliga	female,
visa	see,
uppror	uprising,rebellion,
jul	christmas,
förutsättningarna	prerequisites,conditions,
medan	while,
framgår	will be seen,clear,is shown,
synliga	visible,
våren	spring,the spring,
bred	broad,
bokstaven	the letter,character,
nordöst	north east,northeast,
face	face,
synligt	wisible,seen,visible,
befolkningens	population's,population,
närmade	approached,
brev	letter,
beteende	behaviour,behavior,
uppdelade	divided,
manchester	manchester,
tyvärr	unfortunately,
hopp	hopes,hope,
fursten	prince,
östfronten	eastern front,the east front,eastern,
samisk	samian,sami,lapp,
jan	jan,january,
viktor	viktor,
religionens	religion,religion's,
liksom	and,as is,
jah	jah,
jag	i,
skarsgård	cut farm,skarsgård,
ilska	anger,
handla	act; buy; consume,act,
abba	abba,
parlamentet	the parlament,parliament,
lägger	put,lies,add,
fotbollsspelare	football player,footballers,
lucky	lucky,
generalen	the general,general,
bonde	bonde,farmer,
parlamenten	parliaments,the parliament,
meter	meters,metre,meter,
tidigaste	earliest,
britterna	the brits,british,
h	h,
rowling	rowling,
effekterna	the effects,effects,
iranska	iranian,
rymmer	has,holds,
guvernör	governor,
myndigheterna	authorities,the authorities,the authoroties,
debuterade	debut,debuted,
michail	michail,
konungarike	kingdom,
avlidit	perished,died,
priset	the prize,rate,
kronisk	chronic,
lämplig	suitable,
freddy	freddy,
vietnams	vietnam's,vietnam,
författarskap	the writer,authorship,
sjöng	sang,
upprättandet	establishment,establishing,
tvingade	forced,forcing,
sjönk	sunk,sank,decreased,
balansen	balance,the balance,
varning	warning,
inriktade	oriented,
kategorisvenskar	category swedes,
striden	battle,fight,
finalen	final,
bolivias	bolivia,bolivia's,
strider	strides,conflict,battles,
bilar	car,cars,
ende	only,
förklaringar	explanations,
kedjor	chains,
islamiska	islamic,
ett	a,one; a; an,
marknaden	the market,market,
figuren	the character,figure,
religiöst	religious,
tycker	do,think,thinks,
fåglar	birds,
egypten	egypt,
norge	norway,
etc	etc.,
harvard	harvard,
marknader	markets,
ogillade	disliked,
belägen	located,situated,disposed,
utövade	exerted,exercised,
tätbefolkade	densely populated,populated,
ekvatorn	equator,the equator,
religiösa	religious,
framgången	success,the success,
co	co,
dör	dies,die,
ca	cirka,approximately,
mengele	mengele,
cd	cd,
död	death,dead,dod,
bröllop	brollop,wedding,
stabila	stable,
musikvideo	music video,
cp	cp,
öst	east,
dök	appeared,dove,turned,
antal	number of,number,
jussi	jussi,
keltiska	celtic,
företaget	the company,
moraliskt	morally,moral,
överallt	in all,everywhere,overall; everywhere,
centralort	central city,centralot,regional centre,
växt	plant,
genetik	genetics,
moraliska	moral,
företagen	the companies,taken present,
antas	is required,assumed,expected (to),
antar	adopting,adopt,suppose,
typisk	typical,
frågorna	questions,questions; issues,
molekyler	molecules,
tvungna	forced,forced to,
sänts	sants,sent,
atlanta	atlanta,
friska	healthy,fresh,healty,
haile	haile,
mandatperiod	term,term (of office),term of office,
långsamma	slow,
erhöll	obtained,recieved,acquire,
weber	weber,
rikets	the realms,its,the kingdom's,
demokrati	democracy,
aktivitet	activity,
vd	ceo,
ondskan	the evil,evil,
förlopp	process,pattern,developments,
omnämns	mentioned,is mentioned,
vi	we,
ryssland	russia,
vm	world championship,vm,
lust	desire,loss,
vs	vs,
flickor	girls,
skapare	creator,
föreligger	is,exist,
sitt	his,its,
slovenska	slovenian,
evenemang	event,
spela	play,
tupac	tupac,
armé	poor,army,
känt	known,famous,side,
juan	juan,mr juan,
medeltida	middleaged,medival,medieval,
foundationthe	the foundation,
huden	skin,
paulo	paulo,
matthew	matthew,
und	und,
terrorism	terrorism,
flesta	most,
ball	ball,
columbia	columbia,colombia,
sade	said,
konstantin	konstantin,constantine,
framförde	performed,presented,
nederlag	defeat,
anfield	anfield,
ikea	ikea,
sjukhus	hospital,hospitals,
diabetes	diabetes,
representera	represents,represent,
obamas	obama,obama's,
off	off,
mänskligt	human,
väger	weighs,weight,
vägen	the road,road,
ledde	resulted,led,
ledda	led,run (by),
uno	uno,
versaillesfreden	versailles peace,treaty of versailles,
vägarna	paths,roads (roadways),
gatan	street,the street,
kontakt	plug,contact,
paus	pause,paus,
aktuell	current,
renässansen	the renaissance,renaissance,
paul	paul,
pappa	dad,
tolkade	interpreted,
förknippas	associated to,associated,associate,
kunder	customer,customers,clients,
planeter	planets,
frågan	issue,the question,
englands	england's,
planeten	planet,the planet,
kosovos	kosovo's,kosovo,
filmens	the film's,film,
framtid	future,
förknippad	associated,
motorvägen	motorway,highway,
government	government,
ledarna	the leaders,conductors,
gul	yellow,
dess	then,its,
arbetarklassen	working class,the working class,
tillverkning	production,
pressas	pressed,
följeslagare	companions,companion,
lät	made,had,sounded,
läs	read,
lär	teach,learn,
aktiebolag	companies,limited company; joint-stock company,stock company,
vallhund	herder,herding dog,
stadsbild	cityscape,
amazonas	the amazon rainforest,amazon,amazonas,
symptomen	symptoms,the symptoms,
högskolan	hogs school,university,college,
flotta	fleet,
län	state,between,
tackade	thanked,said/thanked,
bredare	wider,broad,
miniatyr|	miniature,
filmografi	filmography,
anarkismen	the anarkism,anarchism,
trotskij	trotskij,trotsky,
lägsta	lowest,minimum,
stannar	stays,stop,stay,
transport	carriage,transportation,transport,
skriftliga	written,
ockupation	occupation,
februari	february,februari,
kolonin	colony,
behandlades	treated,
toppar	tops,(that) peaks,peak,
sålt	sold,
dags	time,
naturlig	natural,
kollektivtrafik	public transport,
ateist	atheist,
svaga	faint,weak,
fråga	ask,fraga,question,
biologi	biology,
ateism	atheism,
östberlin	east berlin,
svagt	weak,
gandalf	gandalf,
smärta	pain,
vargen	the wolf,
användande	use,use; usage,
kontinenten	the continent,
må	feel,may,mon,
basis	basis,
höger	right,
blodiga	blooded,bloody,
angeles	angeles,
kontinenter	continents,
warner	warner,
solsystemets	solar system,
hittills	date,so far,
burma	burma,
anpassade	adjusted,custom,
släpper	release,releases,
upplösningen	dissolution,disbandment,
sekelskiftet	turn,the turn of the century,
planetens	planet,the planets,
kristus	christ,
lund	grove,lund,
mera	more,
ting	matters,thing,things,
peters	peters,
skola	school,
blå	blue,blah,
fläckar	stain,stains and spots,
bedöms	expected,judged,evaluated,
överbefälhavare	commander-in-chief,supreme commander,
frisk	healthy,fresh,
radioaktiva	radioactive,
samlingar	collections,collection,
förre	pre,former,
uppvisade	showed,
indonesien	indonesia,
apollo	apollo,
socialistiska	socialistic,socialist,
svält	starvation,starvations,
återkommer	will return,returning,
society	society,
official	official,
volvo	volvo,
ruset	the fuddle,intoxication,
stormakt	great power,major power,
monument	monument,monuments,
inrättades	established,were implemented,
problem	problem,problems,
butiker	shops,stores,
ovanför	over,above the,above,
leukemi	leukemia,
heter	units,(is the) name (of),is named,
guy	guy,
utnyttjar	using,uses,
utnyttjas	utilized,used,
skilsmässa	divorce,
separerade	separated,
broder	brother,
banan	the track,banana,
vitryssland	belarus,
månader	months,
sharia	sharia,
programmet	program,the application,the program,
relationer	relations,
distinkta	distinct,
särskilt	in particular,particulary,especially,
relationen	the relation,ratio,
månaden	the month,months,month,
oavgjort	tie,draw,
modernistiska	modernistic,modernist,
bröd	bread,
övergång	transition,
francisco	francisco,fransisco,
uttalade	commented; made a comment; spoke about,spoke,stated,
tider	times; ages,times,
förhandlingar	negotiations,
bröt	brot,broke,
tiden	the time,time,
inspiration	inspiration,
syrgas	oxygen,
syskon	sibling,siblings,
mozart	mozart,
sänker	lowers,lower,sinks,
jordbävning	earthquake,
provinser	provinces,
kommersiell	commercial,
nederländska	netherlands,dutch,
brevet	the letter,letter,
näsan	the nose,nose,
child	child,
elisabeth	elisabeth,
bob	bob,
bosniska	bosnian,
representanthuset	house of representatives,
invadera	invade,
preussen	prussia,
konsekvenserna	impact,consequensis,
smålands	smaland's,småland,
bäst	best,
barmel	barmel,
bibel	bible,insulin,bilble,
spel	game,
edward	edward,
grundande	founding,
ren	deer,clean,
konsekvens	impact,consequence,
mördade	murdered,
konsekvent	consistent,consistency,
grönsaker	vegetables,
golvet	the floor,floor,
främsta	primary; foremost; primarily; principally,request,primary,
främste	chief,premier,
geologi	geology,
jacob	jacob,
skolor	schools,
innefattar	comprises,includes,
uttryck	expression,
upphörde	ceased,expired,discontinued,
estland	estland,estonia,
jamaica	jamaica,
starkast	strongest,
ständerna	the cities,
galax	galaxy,
horn	horns,horn,
colorblack	color black,
alltsedan	even since,since,
förbättringar	improvements,improvement,
eurovision	eurovision,
italiens	italy's,italian,
verksamma	active,
kraftfull	forceful,powerful,
tolv	twelve,
bidrag	contribution,contributions,
nina	nina,
vampyr	vampire,
cyklar	bicycles,bikes,cycles,
bidrar	contributes,
petra	petra,
musikalen	the musical,
räddar	saves,saved,rescues,
bortgång	passing,death,
pluto	pluto,
rapporterar	reports,
norstedt	norstedt,
begått	comitted,committed,
olsson	olsson,
studeras	studied,(is) studied,is studied,
sidan	page,the side,side,
interstellära	interstellar,
regerande	reigning,ruling,
hänvisade	referred,refer,
förblir	remains,remain,
stoft	dust,
träda	esterified,emerge,fallow,
placerades	placed,
akc	akc,
underverk	wonders,wonder,
kongressen	congress,
järnmalm	iron ore,jarnmalm,
fastställdes	confirmed,set,
bro	bridge,
läkemedelsverket	medical products agency,medicines work,food and drug administration,
tillsammans	together,
faktiska	actual,
total	total,
absolution	absolution,
stått	stood,
sarah	sarah,
regenter	monarchs,regents,
negativa	negative,
foster	fetus,fetal,
indiana	indiana,
negativt	negative,
supportrar	supports,supporters,
ifall	if,
förebyggande	preventing,preventive,prevention,
giovanni	giovanni,
fingrar	finger,fingers,
award	award,
riksväg	national highway,highway,
nku	nku,
alces	alces,
inleds	starts,start,
kurderna	kurdish,kurds,
springer	running,springer,
absorberas	absorbed,(gets) absorbed,
friheten	freedom; liberty,freedom,liberty,
beväpnade	armed,
tänkare	thinker,
dokument	files,document,documents,
era	yours,era,
transparency	transparency,
specialiserade	specialized,special,
klorofyll	chlorophyll,cholophyll,
folkmun	popular lore; popularly,common speech,colloquially,
gloria	gloria,
vackra	beautiful,fine,
felaktiga	false,
ekonomiskt	economic,economically,economical,
sommar	summer,
indien	india,
felaktigt	incorrect,erronenous,error,
indier	indians,
enhet	unit,entity,
valborg	may day,valborg,
utlandet	foreign land,abroad,foreign,
gotlands	gotland's,gotland,
solen	the sun,sol,
firas	celebrated,celebrate,
firar	celebrates,celebrate,
gillar	like,enjoy; like,likes,
leonard	leonard,
halland	halland,
beach	beach,
sammansatt	composed,compound,
rädd	scared,afraid,
biografer	movie theaters,movie theaters; cinemas,cinemas,
kategorieuropas	category europe,
lag	law,act,
koreakriget	korean war,the korean war,
visste	did,
tjäna	profit,earn,make,
lat	methacrylate,
law	law,
orden	the words,words,
medlemsstat	member state,
vänsterpartiet	leftist party,left-wing party,left wing party,
lämningar	remains,remnants,
green	green,
massmedia	media,mass media,
livets	life's,life,the life's,
ordet	the word,word,
order	order,
arbetslöshet	unemployment,unemplyment,
natten	overnight,
office	office,
sovjet	soviet,
diagnos	diagnostics,
exempel	example,for example; for instance; sample(-s),
ramadan	ramadan,
söderut	south,
stämmer	(if it's) true,correct,is true,
blandning	mix,mixture,
japan	japan,
bidra	contribute,
vilken	what,which,
straff	penalty,punishment,punishments,
lagets	substrate,the team's,
fragment	fragment,fragments,
vanligtvis	usually,generally,
ämne	substance,
band	band,tape,
fredsbevarande	peace,peacekeeping,
bana	course,web,
they	they,
spelningen	the gig,the concert,
bank	bank,
ansvariga	charge,
huvudartikel	main article,principal article,
l	l,
dåliga	poor,bad,
diskuteras	discussed,is discucssed,
knutpunkt	hub,
tendens	tendency,
dåligt	poor,
område	area,
carlos	carlos,
erbjöd	offered,
germanska	germanic,germanian,
inflytandet	the influence,influence,
koldioxid	carbon dioxide,co,
voddler	voddler,
däggdjur	mammalian,mammal,
rummet	room,
kejserliga	imperially,imperial,
asteroidbältet	asteroid belt,the asteroid belt,
daniel	daniel,
därav	thereof,
trafik	traffic,
bruttonationalprodukt	gross national product,bnp,
oskar	oskar,
vete	wheat,
funktionen	function,the function,
veta	know,out,
sedermera	subsequently,since,
veto	veto,vetoe,
standard	standard,
förmodligen	probably,presumably,
tillbaka	back,
berör	affecting,affect,concerns,
amadeus	amadeus,
ange	set,name,
sprit	liqeur,alcohol,
väldiga	immense,mighty,vast,
professionell	professional,
väldigt	very,
höll	held,hold,gave,
personerna	people; persons,subjects,the persons,
funktioner	functions,features,
önskar	desired,desiring to,wish,
önskan	desired,
another	another,
statskupp	coup,
ingmar	ingmar,
synnerligen	remarkably; particularly,particularly,quite,
drabbade	suffering,affected,
begränsas	limited,(gets) limited,begransas,
begränsar	limit,limits,
ingen	there is no,no,
begränsat	limited,restricted,
sång	song,
förklarade	explained,said,
växthusgaser	vaxthusgaser,greenhouse gas,
inget	not,no,
john	john,
begränsad	restricted,limited,
medborgare	citizens,
antisemitismen	antisemitism,anti-semitism,
äter	eat,eats,
varifrån	from where; wherefrom,from which,
albert	albert,
åland	Åland,
kvarvarande	lasting,remaining,residual,
persson	persson,
bojkott	boycott,
kraftverk	plant,power plant,
trupp	troop,troops,
källkod	source,source code,
militära	military,
religionerna	religions,the religions,
symboliserar	symbolized,symbolizes,
binda	bind,tying,bond,
kronan	kronan,crown,swedish krona,
sonen	the son,
scener	scenes,
används	use,used,
scenen	the stage,stage,
binds	bind,bound,(is) bound,
iron	iron,
byggts	built,
minut	minute,
använde	used,
använda	using,
årens	the year's,years,
skolorna	schools,the schools,
mannen	art,the man,
släktet	the genus,
onani	masturbation,
höja	increase,hoja,raise,
fåglarna	the birds,birds,
omvandling	transformation,
avancerade	advanced,
koloniala	colonial,
anledningar	reasons,
kalendern	calendar,calender,
stavning	spelling,
magnus	magnus,
höjd	height; above,height,
sjukvård	health care,healthcare,care,
aftonbladet	aftonbladet,newsweek,the evening paper,
lades	put,was,
figurerna	figures,characters,
närvaro	attendance,presence,
verkat	worked,acted,seemed,
verkar	acting,seems,operates,
maiden	maiden,
bruce	bruce,
utställning	display,exhibition,
skansen	forecastle,
fjädrar	spring,feathers,
verkan	effect,
flygplatsen	airport,the airport,
aminosyra	amino acid,
vägg	wall,
eviga	eternal,
ägda	owned,
freja	freja,joe,
ägde	tookplace; occured,was,owned,
bortom	beyond,beyond the,
läran	teaching,the teaching,
evigt	forever,eternal,
försvarade	defended,
förväxla	confuse,mistake,
effekten	the effect,effect,
mitten	middle,mid,
damer	ladies,
lewis	lewis,
hinduiska	hindu,
vanligen	usually,typically,
tilläts	was allowed,were allowed to,allowed,
vintrar	winters,
effekter	effects; repercussions,effects,
fortplantning	reproduction,sex,
vätet	hydrogen,the hydrogen,
sättet	manner,way,the way,
 kilometer	kilometer,
sätter	place,puts,sets,
näring	nutrition,
estetiska	aesthetic,
ambassad	embassy,
kejsar	emperor,
inställning	attitude,setting,view,
målvakt	goalee,goalkeeper,
variera	vary,
kontinuerlig	continuous,
imperium	empire,
dj	dj,
di	di,
de	the,they,
dc	d.c.,
sverigedemokraterna	sweden democrats,swedish democracy,
stalins	stalins,stalin,
watson	watson,
människorna	men,the humans,
orolig	worried,
riktningen	direction,denomination,
du	to,you,
dr	doctor,dr,doktor,
sattes	was added,
peyton	peyton,
offret	the victim,offering,
runt	around,between,
emo	emo,
konst	art,srt,
sentida	recent,
splittrades	shattered,split,
offren	victims,
tyngre	heavy,heavier,
fågelarter	bird species,species of bird,
viktigt	important,
libanon	lebanon,
kurdiska	kurdish,
vanlig	ordinary,common,normal,
utförd	completed,performed,
utföra	perform,out,
förena	combine,unite,combining,
väsen	being,entity,
återställa	reset,restore,resett,
präglats	been characterized,been marked,marked,
utfört	done,
massiva	solid,massive,
utförs	out,is done,
sexuell	sexual,
djuret	the animal,animal,
fornnordiska	old nordic,ancient nordic,old norse,
månarna	moons,
fångenskap	captivity,
piratpartiet	pirate party,
djuren	the animals,animals,
materialet	the material,material,
smaken	the flavour,flavor,
osmanska	ottoman,osmanian,ottoman; osmanli,
komplikationer	complications,
we	we,
självständigheten	independance,independence,
intog	seized,occupied,took,
miljö	environment,
jämförelse	comparative,comparison,
huvudsakligen	generally,primarily,
militären	military,the military,
garanterar	ensures,guarantees,
muhammed	muhammed,
kännetecknas	is characterized,characterized (by),characterized,
cox	cox,
kommer	is,
brad	brad,
gruppens	group (-s),group,
målningen	milling,the painting,
samverkan	co,cooperation,
graviditeten	the pregnacy,the pregnancy,
kännetecken	characteristics,distinction,sign,
thierry	thierry,
fångar	captures,prisoners,
tusentals	thousands,
genomför	implement,carry out,out,
tony	tony,
slaveriet	slavery,
smith	smith,
japans	japans,japan's,
patienten	patient,the patient,
biologiska	biological,
lösning	solution,solution; resolution,
framträdande	apperance,appearance,
hitlers	hitlers,
patienter	patients,
klubblag	club teams,club team,
nära	close,near,
attacken	the attack,attack,
vindar	winds,
attacker	attacks,assaults,
fest	festival,party,fest,
juridik	law,
drottningen	queen,the queen,
frekvens	frequency,
bulgariens	bulgaria's,bulgaria,
fromstart	starting from,
vagn	wagon,carrige,
johansson	johansson,
påstådda	said,alleged,
kupp	kupp,coup,coup (d'etat),
aik	aik,
anhängare	followers,supporters,
nordöstra	nordeastern,northeast,
klippa	cut,
release	release,
spanjorerna	spaniards,the spaniards,spanish,
gärdestad	nugent,
have	have,
moldavien	moldova,
deltagarna	the participants,participants,
jordbruk	agricultural,
påverkades	was affected by,affected,
själva	self,actual,
våg	vague,road,wave,
patent	patent,
datorer	pc,
bergskedjor	mountain ranges,
självt	itself,
utgivna	issued,published,
ersattes	was replaced by,replaced,
andelen	share,the share,the proportion,
producerades	produced,was produced,
raid	raid,
hann	did,reached,managed to (in a period of time),
saddam	saddam,
balkan	balkan,the balkans,
sexualitet	sexuality,
delstater	states,
hand	hand,care,
delstaten	land,the state,
nervosa	nervosa,
hans	his,
bilen	the car,car,
koncentrerad	concentrated,concentration,
aspekter	aspects,
förlorade	lost,
rörelsen	movement,
kyla	cold,cooling,
riksdag	parliament; diet,parliament,the parliament,
rör	touch, move(-s),touches,row,
styrkorna	forces,
mamma	mother,
monaco	monaco,
rörelser	movement,movements,
the	the,
röd	red,
thc	thc,
skottland	scotland,
gärningsmannen	perpetrator; offender,the offender,culprit,
newton	newton,
kall	cold,
nästan	almost,close,
kroppens	the body's,the bodies,
goda	good,
enades	agreed,
kalender	calendar,calender,
upptäckte	discovered,found,
swahili	swahili,swahilli,
lindh	lindh,
så	as,so,
distributioner	distributions,
snus	snuff,
wright	wright,
havets	the seas,sea,
skick	state,condition,
kvinnan	woman,female,
samfund	communities,order,
plasma	plasma,
viking	viking,
förbättra	improve,
föda	feed,give birth; food,give birth,
återgick	returned,returning,
skadorna	injuries,damages,damage,
arab	arab,
fusion	fusion,
indianer	indians,
föds	born,
everton	everton,
picasso	picasso,
hepatit	hepatite,hepatitis,heptatitis,
acceptera	acceptable,accept,
årlig	yearly,
indelning	the subdivision,classification,
indelningen	division,subdivision,classification,
dahlén	dahlén,
xbox	xbox,
gandhi	gandhi,
transkription	transcription,transcript,transcripton,
sixx	sixx,
motsvarighet	equivalent,
avsätta	unseat,depositing,
bort	away,remove,
born	born,
presidentvalet	presidential elections,presidential election,
borg	tower,castle,
bord	table,
kungar	kings,
humor	humor,humour,
territorierna	territories,
purple	purple,
serbiens	serbias,
siffran	figure,the number,number,
vinterkriget	the winter war,winter,winter war,
columbus	columbus,
stadsdelarna	districts,neighborhood (-s),
vägar	roads,paths,
trosbekännelsen	creed,faith of confession,
fängslades	imprisoned; jailed, gaoled; incarcerated,jailed,
post	week,not a swedish word,
slovakien	slovakia,
vunnit	win,won,
upplösning	resolution; dissolution,resolution,
banker	banks,
olika	different,variety,
jacques	jacques,
återfinns	found,is rediscovered,
samer	sami,
roms	romes,roms,rome's,
lois	lois,
epicentrum	epicentre,epicenter,
kommittén	the committee,committee,
blivande	prospective,future,to be,
gemenskapen	the collective,community,
way	way,väg,
was	was,
war	war,
representerar	represents,
hypotes	hypothesized,hypothesis,
skiljas	separated,separate,
motorvägar	highways,motor,
inträffar	occurs,occur,
inträffat	occurred,
partiledare	party leader,
emil	emil,
reser	travels,rise,rises,
studierna	studies,the studies,
mtv	mtv,
finansiering	financing,financiation,
litterär	literary,
långvarig	of long duration,prolonged; lengthy; long,long,
träning	training,practice,
erövra	conquer,
engagerade	dedicated,engaged,committed,
moore	moore,
utomlands	abroad,
tesla	tesla,
xiis	xii,
efter	after,
bilderna	the pictures,
xiii	xiii,
moln	cloudy,cloud,
empati	empathy,
toppen	top,peak,the top,
alltid	always,
möta	meet,face,
förmåga	abilities,ability,
janukovytj	janukovytj,yanukovych,
möte	meeting,
arkitekter	architects,
test	test,
götaland	götaland,gotaland,
konservatism	conservatism,
mött	faced,met,
femton	fifteen,
tottenham	tottenham,
räknat	calculated,counted,
reglerar	regulates,controls,
regleras	controlled,regulated,is regulated,
rätter	dishes,
hemma	home,at home,
omgivande	surrounding,surounding,ambient,
rätten	right,the court,
solens	the sun,solar,
bergmans	bergman's,bergmans,
dance	dance,
uppfanns	was invented,invented,
tenderar	tend,
datum	date,
förklaringen	the explanation,statement,
osäker	insecure,unsure,
lider	suffering,suffers,
utkämpades	fought,
förhistorisk	forhistorisk,prehistorian,
afrikaner	africans,
heller	neither,neither; nor,nor,
rådet	the council,council,
igelkott	hedgehog,
zone	zone,
vattenånga	steam,water vapour,
ätten	the dynasty,dynasty,
terror	terror,
vänder	turn,face,
brown	brown,
charles	charles,
hannah	hannah,
uttrycka	express,
enskild	single,
lättare	light,easier,
hannar	males,
vegas	vegas,
uttryckt	expressed,
avbröts	canceled,interrupted,
enskilt	individually,single,
salvador	salvador,
stycken	pieces; parts,pieces,
gud	god,
nedsatt	impaired,reduced,decreased; diminished,
datorspel	video game,computer game,
hisingen	hisingen,
levnadsstandard	living standard,standard of living,
frigörs	released,is released,
ljuset	the light,light,
säte	sate,seat,
formella	formal,
litterära	literary,literal,
templet	the temple,temple,
revolution	revolution,
alfa	alpha,
cosa	cosa,
engagerad	dedicated,engaged,
invandrade	immigrated,immigrant,
sköttes	operated,handled,
mål	case,goal,mal,
formellt	formally,formal,
motsatte	opposed,
midsommar	midsummer,
stimulera	stimulate,stimulating,
motsatta	opposite,
yorks	yorks,
ungdomar	youths,adolescents,the youth,
tidig	early,
ingick	were included,was,
kosmiska	the cosmic,cosmic,
uniform	uniform,
fastigheter	real estates,properties,
utspelar	takes place,set,
versionen	edition,the version,
gener	genes,
muslim	muslim,
marxismen	marxism,the marxism,
kärlek	love,
påstås	claimed,(been) said,allegedly,
klassificeras	classified,
genen	gene,the gene,
oerhört	tremendously,extremely,
tillträde	access,
antarktiska	antarctic,
flames	flames,
sistnämnda	later,last,
kemi	chemistry,
franklin	franklin,
ponny	pony,
fronten	front,the front,
vinnare	win,winner,
ekr	ekr,ad,
churchill	churchill,
marken	soil,
extra	optional,extra,
vapnet	the weapon,the weapon; escutheon; coat of arms; arms; badge,
spridit	spread,disseminated,
konkret	specific,concrete,
ukrainas	ukranian,ukraine's,ukrainian,
vapnen	weapons,the weapons,
förteckning	index,listing,label,
fbi	fbi,
kärnkraftverk	nuclear power plant,nuclear powerplant,
presenterar	presents,present,
upprättade	established,prepared,
äktenskapet	marriage,
super	super,
territorier	territories,
stabilitet	stability,
live	live,
regel	rule,
territoriet	territory,
angels	angels,
överhuvudtaget	on the whole,in general,in general, generally,
fransmännen	the french,frenchman,french,
parallellt	at the same time,parallel,
club	club,
rivalitet	rivality,rivalry,
snabbt	fast,quickly,
enda	only,single,
målvakten	the goalkeeper,
zarathustra	zarathustra,
ämnena	subjects,the elements,substances,
närmar	close,closing,close in,
varför	therefore,why,
kolonialismen	the colonialism,colonialism,
feministiska	feminist,
snabba	rapid,fast,
löner	wages and salaries,salaries,
ibm	ibm,
ibn	ibn,
interaktion	the interaction,interaction,
frukt	fruit,fruits,
can	can,cancer,
erbjuder	offers,
heart	heart,
några	few,a few,
december	december,
nobels	nobel,nobel's,
influensavirus	flu virus,influenza,flue virus,
gentemot	towards,against,
abort	abortion,
uppstår	occur,
genomgått	experienced,passed,
ligan	league,
pojke	boy,
uppskattades	estimated,appreciated,was appreciated,
betydelse	importance,significance,
kopplingar	connections,links,
perserna	the persians,persians,
southern	southern,
riktlinjer	guidelines,
framgångarna	successes,the successes,
göteborgs	gothenburg,gothenburgs,
gräns	limit,border,
ungern	hungary,hungaria,
förutsättning	provided,prerequisite,
romarna	romans,the roman,the romans,
flyttas	is moved,moved,
flyttar	move,
kurt	kurt,
kurs	course,rate,
michel	michel,
ukrainska	ukrainian,
rekordet	record,the record,
maktens	the powers,forces,the power's,
landshövding	county governor,governor,govenror,
ingripa	interfere,act,
ganska	rather,fairly,quite,
ättlingar	descendants,
magnetfält	magnetic,magnetic field,
generalguvernören	governor-general,governor general,general governor,
linnés	linnaeus,
fält	field,
skabb	mites,scab,scabies,
idéerna	ideema,ideas,
levde	lived,survived,
utnämndes	was declared,appointed,
därifrån	from thence,from there,
bergskedjan	mountain range,the mountain group,
nominerades	was nominated,nominated,
hals	throat,neck,
varav	of which,which,
arton	18,eighteen,
halv	half,
nog	sufficiently,enough,
författarna	the authors,writers,
förvaras	stored,is stored,
komponenter	components,
begränsa	limit,
not	note,
nou	nou,
rakt	straight,
now	now,
dödsstraffet	capital punishment; death penalty,death penalty,the death penalty,
hall	hall,
frihet	freedom,
james	james,
språk	language,
främmande	foreign; alien,undesirable,foreign,
antyder	indicates,
stockholm	stockholm,stocholm,
januari	january,
drog	draw,pulled,drug,
aspergers	downs syndrome,aspergers,
em	em,european championship,
el	el,
en	a,
flamländska	flemish,
ej	not,no,
ed	ed,
eg	ec,
utbrett	wide,widespread,
spåra	track,trace,
strålningen	the radiation,radiation,
ex	eg,ex,
kroatiska	croatian,
et	et,
resultera	result,
fuglesang	fuglesang,
ep	ep,
premiärministern	the prime minister,prime minister,
er	you,your,
album	album,
teorier	theories,
återkommande	recurring,
hustrun	the wife,his wife,
kortare	shorter,
stallone	stallone,
punkt	item,point,
genetisk	genetic,
taget	a time (practically; virtually; any; at all),time,
välkänd	known,well-known,well known,
marina	marina,marine,
betraktades	considered,regarded,
böhmen	bohemia,
british	british,
domen	judgment,verdict; judgement,
linné	linen,linneus,temperature,
fc	fc,
allmänheten	public,general public,
arbetsgivare	employers,
skådespelerska	actress,
xi	xi,
förändrats	changed,
derivatan	derivative,the derivative,
ring	ring,
xv	xv,
bergqvist	bergqvist,
våglängder	wavelength,wave lengths,wavelengths,
omtvistat	contentious,disputed,controversial,
priser	rates,prizes,
desmond	desmond,
svenske	swedish,
sheen	sheen,
dessutom	moreover,furthermore; moreover, additionally; likewise,furthermore,
satsningar	ventures,investments,resources,
färre	fewer,less,
that	that,
nödvändig	necessary,essential,
fascisterna	the fascists,the facists,fascists,
delats	divided,been awarded,
television	television,
europeisk	european,
sidorna	the pages,pages,
utbyggda	expanded,expand,
ändrades	changed,was,
yttre	outer,
grundad	founded,based,
craig	craig,
premier	premiums,
statsminister	prime minister,
faktor	factor,
kairo	cairo,
grundat	founded,(was) found,based,
grundar	bases,based,
grundas	is based,based,
anger	indicates,gives,
anges	mention,is put at,specified,
befolkningstillväxt	population growth,befolkningstillvaxt,
hjälp	using,help,
hör	include,belong,hears,
själv	alone,own,himself,
skär	will,cut,skerry,
fortsatte	continued,
fortsatta	continued,
etiopiska	ethiopian,etiopian,
bönor	beans,
hög	high,
online	online,
skäl	reasons,reason,
kategoriorter	category visited,
numera	now,nowadays,
santiago	santiago,
successivt	successively,progressively,
egentlig	actual; factual; real,actual,
bekostnad	detriment,expense,
dvärgar	dwarves,dwarfs,
glödlampor	lightbulbs,light bulbs,filament,
america	america,
på	on,in, on, at,
michelle	michelle,
lyfter	lift,lifts,lifting,
norrmän	norwegians,
nordligaste	northermost,northern,northernmost,
parlamentets	the parliament's,parliament,
runda	round,
orsaka	cause,
abraham	abraham,
skapats	was created,generated,
doktor	doctor,
kyrkorna	churches,the churches,
nazisternas	the nazi's,nazi,
marocko	morocco,marocco,
colombo	colombo,
teori	theory,
perfekt	perfect,
mannens	man,man's,
byggda	constructed,
rötter	roots,
varmblod	warmblood,warm-blooded,
adolf	adolf,
raúl	raul,
himmel	heaven,
huskvarna	huskvarna,
epoken	epoch,the epoch,
dagbok	diary,log,
sierra	sierra,
mörk	dark,
definierade	defined,
uppståndelse	resurrection,
helgdagar	holidays,
riddare	knight,
samuel	samuel,
gudarnas	the gods',gods,god's,
ambitioner	ambitions,
folkomröstning	referendum,
marxistisk	marxist,marxistic,
tävla	compete,
handlingar	actions,
drabbas	troubled with,suffer,affected,
facupen	fa cup,fa-cup,
längst	at,farthest,longest,
bushadministrationen	the bushadministration,the bush administration,bush administration,
länge	long,
storstäder	metropolises,cities,
kommande	upcoming,
tillfällig	temporarily,
osbourne	osbourne,
övergången	transition,the transition,transformation,
sport	athletics,sport,
katastrofer	disasters,catastrophes,
depressionen	the depression,depression,
konstaterade	concluded,established,stated,
ladin	ladin,
depressioner	recessions,depressions,depression,
israels	israels,israeli,israel's,
import	import,
kommunismens	communism,the communisms,the communism's,
katastrofen	catastrophy,the catastrophy,disaster,
yta	surface,
ronja	ronja,
personlighet	character,personality,
flygande	flying,
männen	the men,men,
utgivningen	release,the publication,the release,
verket	plant; indeed,plant,board,
hendrix	hendrix,
verken	plants,wroks,
utgavs	was published,published,
comeback	comeback,
samtal	conersation,call,
monicas	monica,monica's,
mona	mona,
bördiga	fertile,
placerad	placed,disposed,
handlar	is,concerns,
kristinas	kristina's,crisis thawed,
propaganda	propaganda,
feminismen	feminism,
ståndpunkt	standpoint,position,
nils	nils,
comet	comet,
placerar	place,places,
placeras	placed,
utnyttja	use,
avskaffande	elimination,abolition,abolishment,
dömande	sentencing,judging,
regeringens	government,government's,
lägenhet	apartment,appartment,
bomull	cotton,
riksrådet	riskradet,privy council; council of state; crown council; senate,privy council,
östtyska	east german,
överlever	survives,
handlande	action,
långfilm	feature film,feature movie,
oliver	olives,
välstånd	prosperity,
wien	vienna,
karlstads	karlstad's,
sker	happens,is,
oden	node,oden,
knappt	barely,
försörjde	living,provided,
dräkt	costume,outfit,
observera	note,observe,
utförda	formed,performed,made,
riktningar	directions,direction,direction (-s),
elvis	elvis,
funnits	found,been,
ik	ik,
konservativa	conservative,
ytan	the area,surface,area,
uefacupen	the uefa champions league,uefa europa league,uefacupen,
rapporter	reports,
prinsessan	the princess,princess,
rapporten	report,the report,
polens	polands,pole,
ordningen	the order,order,procedure,
ändå	still,spirit,
ansikte	face,
tjeckien	czech republic,the czech republic,
eran	era,
beläget	located,base,
inslag	impact,elements,element,
finanskrisen	financial crisis,the financial crisis,
tänkande	thinking,
behandlade	was treated,treated,
kvarter	quarter,block,neighborhoods,
kenya	kenya,
västerländska	vasterlandska,western,
katalanska	catalan,
helium	helium,
grundade	founded,based,
infödda	natives,native,
slaget	the strike,type,
långt	far,long,
orsakade	caused,causing,
programvara	software,
media	media,
långa	langa,long,
talmannen	president,speaker of the riksdag,
homosexualitet	homosexuality,homosexuallity,
kromosom	chromosome,
pesten	the plague,death,plague,
lite	little,a little,
figurer	figures,
speciella	special,
offensiven	offensive,the offensive,
begär	requests,request,
skivbolaget	record label,the record company,
acdc	ac/dc,
omfattande	wide-ranging,large,massive; extensive,
målningar	paintings,
omfattas	comprise,subject,
speciellt	particularly,
omgående	immediately,immediate,
ekonomisk	economic,
tradition	tradition,
fredspris	peace prize,
skånes	scania,scania's,
erkänd	acknowledged,recognized,
erkänt	recognized,
flaggor	flags,
kategorilevande	category of live,
mynning	outfall,muzzle,mouth,
forskarna	the scientists,scientists,
skandinaviska	scandinavic,scandinavian,
tydlig	clear,obvious,
botten	the base,bottom,
samiska	sami,
eleverna	the pupils,the students,
lagerkvist	lagerkvist,
spänningar	tensions,
nazismen	nazism,
euron	the euro,euro,
malcolm	malcolm,
lade	laid,added,seized,
ditt	your,
strävar	striving; aiming (to; for),strives,
irland	irland,ireland,
arbeta	work,working,
stund	while,momentum,
östergötland	Östergötland,east gothland,
selma	selma,
amy	amy,
lady	lady,
tobak	tobacco,
strävan	will,the quest,endeavor,
nationella	national,
skilda	seperated,separate,
miniatyr|en	thumbnail,a minature,
skilde	divided,varied,there was a separation,
varandra	each other,
nationellt	national,nationally,
t	t,e.g.,
låga	cook,low,
astronomer	astronomers,astronomer,
lågt	low,
präglades	was marked,imprinted,marked,
stånd	in the context: (make) the war happen,position,
fönster	windows,window,
slår	states,switch,beats,
användbara	usable,useful,
sålts	sold,
indikerar	indicates,
frigörelse	liberation,
berodde	was,depended,depended upon,
innebörden	meaning,the significance,
bestämd	fixed,
strindberg	strindberg,
utskott	committee,organ,
bestämt	decided,particularly,
nsdap	nsdap,
inuti	inside,
växa	growth,grow,wax,
kategoriledamöter	category members,category: members,
bestäms	determined,is decided,
kaffet	coffee,the coffee,
francis	francis,
övertygad	confident,
ideologi	ideology,
jamaicanska	jamaican,
central	central,center,
bidraget	contribution,grant,
sri	sri,
torget	square,the square,torget,
bidragen	the contributions,contributions,
efterkrigstiden	the post-war period,post-war era,post-war,
kapten	captain,
klassiker	classics,classic,
transporter	carriage,transports,
karriär	career,
your	your,
fast	solid,though; although; fixed; permanent,even though,
area	area,
satsade	invested,bet,
sats	theorem,kit,
stark	strong,
start	start,
anställd	employed,hired,
specifika	specific,
likväl	nevertheless,still,as well,
gånger	times,
fastställa	determine,confirm,
hawking	hawking,
guillou	guillou,
wailers	wailers,
sämsta	worst,
gången	time,
traditionerna	traditions,the traditions,
expeditionen	the expidition,expedition,
spänner	spanner,span,
minne	memory,
engelskan	the english,english,
indelningar	divisions,classifications,
minns	remembers,remember,
miguel	miguel,
bilmärke	car make,make of car,
expeditioner	expeditions,
kostar	costs,
kungen	king,the king,
grammis	grammy,
sveriges	swedens,sweden,
godkände	approved,
styrde	steered,
knut	knut,knot,
transportera	transport,
nere	down,low,
mongoliet	mongolia,
efteråt	afterwards,
upphovsman	creator,author,
tänderna	teeh,teeth,
you	you,
köper	making,
knä	knee,knees,
drift	operation,drift,
översätts	translated,translate,is translated,
massachusetts	massachusetts,massachussetts,
röda	red,
bandmedlemmarna	band members,have,
riktat	directed,pointed,
tjänare	servant,
handelsmän	merchants,
morgonen	the morning,am,
färdas	travels,
susan	susan,
olympiastadion	olympa stadium,olympic stadium,
monte	assembly,
eriksson	eriksson,
beskrivningar	description,descriptions,
energikälla	source,energy source,energy call,
messi	messi,
öknen	the desert,desert,
loppet	bore,the race,
antoinette	antoinette,
griffin	griffin,
råvaror	raw,wood,raw materials,
lämpliga	suitable,
påbörjades	commenced; begun,initiated,was started,
lämpligt	suitable,
fästning	fortress,
skiljer	differs,is different; differ,different,
vers	verse,
jensen	jensen,
får	may be,can,allow,
verk	work,works,
osv	etc.,
spår	track,pairs,
heaven	heaven,
sverige	sweden,
behöver	need,
louis	louis,
manager	manager,
industrialiseringen	indutrialization,industrialization,
resan	the trip,journey,
rasism	racism,
magdalena	magdalena,
skiva	record,disc,
fåglarnas	the birds',birds,
egendom	property,
kritiserats	criticized,critized,
orgasm	orgasm,
markerade	selected,marked,
trupper	troops,
utåt	outwardly,out,
pythagoras	pythagoras,
tvskådespelare	tv actor,
besöker	visit,visits,
bedrev	conducted,managed,
fjärde	fourth,
förbjuden	smoking,
bernhard	bernhard,
förbjuder	prohibiting,forbids,
misstänkta	suspected,suspect,
inblandad	mixed,
förbjudet	prohibited,
irak	iraq,
ersatt	replaced,
iran	iran,
genomförde	carried out,
ersättare	alternate,replacement,
kronor	kronor,crowns,
observeras	observed,is noticed,is observed,
ontario	ontario,
uttalat	pronounced,outspoken,expressed,
lämna	leave,supply,
uttalas	pronounced,be pronounced,
arena	arena,
medarbetare	employees,coworker,
signifikant	significant,
vår	spring,
krigen	the wars,wars,
dyker	dives,shows,
stulna	stolen,
minst	at least,
boxning	boxing,boxing; pugilism,
sagor	fairytales,tales,fairy tales,
kriget	the war,war,
hoppades	hoped,
perspektiv	perspective,
medicin	medicine,
då	then,when,
globen	lobe,the globe,
nazityskland	nazi germany,
gick	went,passed,
grunda	found,base,
dalarna	valleys,dalarna,
ökat	increased,
nukleotider	nucleotides,nucleotide,
familj	family,
avsedd	adapted,intended,
avgör	decides,determines,
simba	simba,pool,
arrangemang	arrangement,
taket	the roof,ceiling,
tillät	distillate,allowed,
etablerad	established,
förlängningen	elongation,
planen	the field,the plan,plan,
trummisen	the drummer,drummer,
oecd	oecd,
bolagets	company's,the corporation's,
representeras	represented,
expansionen	expansion,the expansion,
teatrar	theaters,
massan	mass,
kurdistan	kurdistan,
reptiler	reptiles,
okänt	unknown,
utökat	extended,expanded,
blodtryck	blood pressure,
ständiga	permanent,constant,
latinamerikanska	latin-american,latin american,
site	site,
inspelad	recorded,
räknar	counts,counter,
räknas	calculated,counted,are counted,
lagstiftande	legislative,legislating,legislation,
ständigt	always,constant,
mördad	murdered,murderd,
företeelser	phenomena,
gazaremsan	gaza strip,the gaza strip,
ombord	onboard,board,
livslängd	life,life expectancy,
istället	instead,instead of,
rapporterade	reported,
kejsardömet	empire,
partner	partner,
herrens	lord,
species	species,
zanzibar	zanzibar,
ökar	increases,
gälla	valid,be valid,
serber	serbs,
ledger	ledger,
linköping	linköping,
smitta	infection,
reidars	reidars,reidar's,
ytterligare	further,additional,
samarbetet	co,cooperation,the collaboration,
utför	perform,out,
turkarna	turks,the turks,
torde	could,should,
fastän	although,
försök	experiments,expirements,
utom	except,out,
fd	former,ex,
ff	ff,
invasion	invasions,invasion,
samarbeten	cooperations,collaborations,
fn	un,the un,fn,
stabil	stable,
vattenkraft	water power,hydroelectric power,hydro,
kostnaden	cost,
byggandet	construction,the building,
skivan	record,the record,disc,
enzymer	enzymes,
allmänna	general,
korset	cross,
kognitiv	cognitive,
segrar	wins,victories,
skiljs	separated,separate,
kostnader	cost,expenses,costs,
dream	dream,
nämnts	mentioned,above,
tillgångar	assets,
helt	completely,totally,
bloggar	blogs,
tornet	tower,the tower,
tornen	towers,the tower,
hela	entire,full,
maffian	mafia,
hell	hell,
skillnaderna	the differences,differences,
eros	eros,
hundratusentals	hundreds of thousands of,hundreds of thousands,
romance	romance,
kompositörer	composers,compositors,
antagits	adoption,adopted,
systems	systems,system,
österrikes	austria's,austrias,
mahatma	mahatma,
musikalisk	musical,
bytte	changed,changed it's,swapped,
elden	fire,the fire,
lyckas	successful,succeed,
konstitutionella	constitutional,
greps	was arrested,arrested,(was) arrested,
dyrt	a high price,expensive,dearly,
petter	petter,
närmare	further,close to,
fullt	full; fully; completely,completely,full,
fulla	full,complete,
skrivit	written,wrote,
strålning	radiation,
kontinentens	the continents,continent,
ifk	ifk,
etnisk	ethnic,
neil	neil,
positionen	position,the position,
märktes	labeled,
noga	carefully,
positioner	positions,
rättvisa	justice,
försäljning	sales,sale,
aktörer	players,actors,
robert	robert,
bodde	lived,
lungorna	lungs,the lungs,
stödet	support,the support,
stöder	supporting,supports,
känna	known,know,
utredningen	investigation,the investigation,
heroin	heroin,heroine,
känns	feels,felt,
delningen	division,pitch,
vasas	vasa,vasas,vasa's,
svarade	answered,said,accounted (for); answered,
åtskilliga	several,
etnicitet	ethnicity,ethnic,
skogen	woods,forest,
skilja	seperate,differ; differentiate,separate,
american	american,
förbättrade	improved,improve,
underhåll	support,entertainment,allowance,
kung	king,
sänder	broadcast,transmits,
sändes	was sent,sent,
utvecklats	developed,
synen	the view,sight,
etiska	ehtical,codes,
arsenal	arsenal,
riksföreståndare	regent,
minoritetsspråk	minority language,minority,
fabriker	plants,factories,
helsingborgs	helsing borg,helsingborg's,
taggar	spikes,tags,thorn, twig,
synes	seems to,apparently,appears,
miss	miss,
rygg	back,backs,dorsal,
deltagare	contestant,participants,participiant,
kanada	canada,
kongresspartiet	congress party,indian national congress,
station	station,
parlamentsvalet	parliament election,election to parliament,parliamentary elections,
nigeria	nigeria,
brittiska	british,
luminositet	luminosity,
brittiske	british,
åkte	went,relegated,
lupus	lupus,
förnuftet	reason,the common sense,
brittiskt	brittish,british,
tvungen	forced,had,forced (to),
bildande	forming,founding,formation,
växterna	plants,
stora	large,big,
långsamt	slowly,
aristokratin	the aristocraty,aristocracy,
andersson	andersson,
värden	values,
värdet	the value,
stiftelsen	foundation,
gren	crotch,branch,
sekunder	seconds,second,
charlotte	charlotte,
bestämdes	was decided,decided,was determined,
teslas	teslas,tesla's,
genomgripande	radical,good,comprehensive; radical,
medeltemperaturen	median temperature,the average temperature,
tvärtom	on the contrary,contrary to,vice versa,
nominerad	nominate,nominated,
militär	military,
karl	karl,
vädret	weather,the weather,
grundarna	founders,
liberalismen	the liberalism,liberalism,
henne	she,her,
liv	life,
mänskliga	human,
herre	lord,master; lord,
avseenden	respects,regard,
jämföras	comparable,compared,
mexiko	mexico,
logotyp	logo,logotype,
sektor	sector,
säsongens	season,the seasons,
kan	can be,
bistånd	aid,assistance,
kap	chapter,cape,
fågel	bird,
utgör	make up,constitutes,
himlakroppar	celestial bodies,
södra	southern,south,
läst	read,load,
polacker	polish,poles,
klädd	clothed,coated,
räknade	calculated,counted,
recensioner	reviews,
rådde	prevailed,was,
två	two,
osäkra	insecure,uncertain,doubtful,
ingenting	nothing,
jupiters	jupiter's,jupiter,
möjligen	possibly,
counterstrike	counterstrike,
hänvisar	reference,
muslimsk	muslim,muslim; muslem,
integritet	integrity,
sanna	true,
justice	justice,
humanistiska	humane,humanistic,humanist,
åländska	Åland swedish,aland,
ikon	icon,
lennon	lennon,
darwin	darwin,
ingå	be a part,include,be included in,
dominans	dominant,dominance,
arabvärlden	the arab world,arab world,
tillhört	belonged,belonged to,
utrikes	foreign,
gått	gone,passed,
alexander	alexander,
dogs	dogs,
restauranger	restaurant,restaurants,
avsaknaden	absence,
dömdes	sentenced,was convicted,
vilket	which,
målare	grinders,painter,
x	x,
tolkiens	tolkien,tolkien's,
västkusten	the west coast,west coast,
grunden	base,basis,
allmänt	generally,generally; public,commonly,
maurice	maurice,
ansvar	responsibilities,responsibility,
bakgrund	bakground,background,
tidigare	earlier,before,
ändamål	object,purpose,
grunder	bases,
mörkare	darkey,darker,
förekom	was,
flyter	float,flows,
direktör	director,
haddock	haddock,
pictures	pictures,
lösa	solve,
pjäser	checkers,plays,
löst	solved,dissolved,1st sentence: loosely; 2nd & 3rd: solved,
produkten	product,the result,
chansen	chances,chance,
kategorin	category,the category,
allvar	earnest,serious,
likhet	similar,resemblance,like,
utsträckning	extent,
köket	cuisine,the kitchen,
genre	genre,
länk	link,
produkter	products,
league	league,
lejonet	the lion,lion,
anor	ancestry,lineage; ancestry,
viljan	will,te will,
slavar	slaves,
kyrkliga	religious,from the church,church,
bott	lived,lived in,
läsaren	the reader,reader,
evolutionsteorin	theory of evolution,
uppfylla	satisfy,fulfill,meet (requirements),
betydde	meant,ment,
derivata	derivative,
scientologikyrkan	the church of scientology,church of scientology,
linux	linux,
sokrates	socrates,sokrates,
nacional	nacional,
skydd	protection,
händerna	the hands,hands,
merparten	most,the majority,larger part,
minskade	minimum period,was reduced,
enheten	the unit,unit,
enheter	units,
kuster	coasts,
konsensus	consensus,
gestalt	character,figure,
walter	walter,
isolerade	isolated,
handlingen	hand-writing,the plot,the story,
budgeten	budget,the budget,
anthony	anthony,
livet	the life,life,
delades	shared,divided,split,
genomförs	implemented, carried through,conducted,is carried out,
socialism	socialism,
belgrad	belgrade,
hegel	hegel,
läses	read,is read,
läser	read,are reading,
diktator	dictator,
mängden	amount,the amount,
tillfället	to the case,time,
slutar	ends,end,
slutat	ended,left,
uttryckte	expressed,
nationalitet	nationality,
klippiga	rocky,
sorter	kinds,varieties,types,
bärande	wearing,leading,fundamental; wearing; supportive,
lagar	laws,
tillfällen	occasion,oppertunities,jobs,
kombineras	combined,
staffan	staffan,
kombinerat	combined,
grant	word,
borgerliga	bourgeois,conservative,
deltagande	participation,
sammanlagt	a total of,total,totaly,
nöd	distress,emergency,
demokratin	the democracy,democracy,
kombinerad	combined,
grand	grand,
ingår	is,penetrations,
luxemburg	luxembourg,luxemburg,
folkslag	kind of people,peoples,
kungahuset	royal family,royal house,
bon	nests,bon,
anklagats	accused,
 km	kilometers,
kommunicera	communicate,communicating,
förlag	publishers,magazine,
seglade	sailed,
armenien	armenien,armenian,armenia,
svealand	svealand,
fatta	make,to make,
kurdisk	kurdish,
stjärnorna	stars,the stars,
präglas	characterised,characterized,
cruz	cruz,
frihetliga	libertarian,
flygplan	aircraft,airplane,
nutid	present day,present,
präglad	characterize,marked,characterized,
följande	following,the following,
feminister	feminists,
hotell	hotel,
njurarna	the kidneys,kidney,
tortyr	torture,
skal	shell,skin,
fredliga	peacefull,peaceful,
inlett	started,ushered in,
uppfinnare	inventor,
kallblod	cold blood,cold blooded,draught horse,
taiwan	taiwan,
lik	similar,alike,
gänget	the group,the gang,gang,
nikki	nikki,
barack	barack,barracks,
välkända	known,well known,
varuhus	warehouse,department store,
egenskap	trait,ability,seeks,
djup	deep,
marco	marco,
bestå	consists,exist,comprise,
lika	similar,alike,equal,
gör	does,makes,
kulturen	culture,the culture,
enklare	easier,simpler,
kulturer	cultures,
gitarristen	the guitarist,guitarists,
game	game,
baserade	based,
unga	young,
emma	emaa,emma,
immigranter	immigrants,
innan	before,
uppvärmningen	the warmup,heating,the warm-up,
känslig	susceptible,
releasedatum	release date,
dylikt	such,
koden	the code,code,
infektion	infection,
criss	criss,
gandhis	gandhi's,gandhi,
terminologi	terminology,
unge	young,kid,
history	history,
donna	donna,
begärde	called,demanded,
tolkats	interpretation,interpret,interpreted,
kommenterade	comment,commented,
byggnader	buildings,structures,
biträdande	assistant,assisting,deputy,
pierre	pierre,
våldet	the violence,violence,
economic	economic,ecomomic,
publiceringen	the publication,publishing,publication,
syndrom	syndrome,syndrom,
sammanhängande	context of,connective,continous,
skapat	created,
världsarvslista	world heritage list,
vilda	wild,
skapar	creates,
skapas	creates,
faktorn	factor,
slash	slash,
skapad	created,
enormt	gigantic,fusionenormously,
bägge	both,
sarajevo	sarajevo,
run	run,
steg	rose,step,
rum	(took) place,room,
sten	stone,
mellankrigstiden	interwar years,time between the wars,interwar period,
naturvetenskapliga	science,scientific,
offside	offside,
skrivet	written,
benfica	benfica,
freddie	freddie,
führer	fuhrer,fuehrer,
förtroende	confidence,trust,
myndighet	authoroty,authority,
övergick	transended,went over,switched,
linjen	the line,line,
etablerade	established,
fysiologiska	physiological,
efterträdare	successor,
refererar	refer (to),references,reference,
linjer	routes,lines,
edvard	edvard,edward,
länderna	states,the countries,
ändringar	edit,starts to process,changes,
ida	ida,
fåtal	few,a few,
stanna	stop,stay,
egenskaper	characteristics,charactiristics,qualities,
ön	island,the island,
öl	beer,
reaktorer	reactors,
semifinalen	the semi-final,semi finals,semifinal,
institut	institute,institution,
emellan	a,inbetween; between,between,
överst	top,at the top; uppermost,
föreningen	the association,association,compound,
fokuserade	concentrated,focused,
ligga	lies, lie,lie,be,
spänningen	exitement,voltage,
visas	is showed,shown,
visat	found,shown,
heritage	heritage,
spridd	wide spread,widespread,spread,
jonsson	jonsson,
orsaker	causes,
ledamot	member,representative,
strukturen	the structure,structure,
japanerna	japanese,the japanese,
spektrumet	spectrum,
larry	larry,
strukturer	structures,structure,
drabbats	affected,afflicted,
skådespelaren	actor,
skull	sake,
ute	absent,out,
nyval	re-election,new election,election,
skuld	liability,debt,guilt,
malin	maleic,malin,
trafikerade	traffic,frequent,trafficked,
  km²	square kilometre,km²,km2,
politik	politics,policies,
förbjöds	banned,forbidden,
chelsea	chelsea,
ligacupen	league cup,
bränslen	fuel,fuels,
ihåg	remember,
avsåg	meant,intended,mean,
voltaires	voltaire,
uppfyller	fulfills,
hårdrock	hard rock,hardrock,
igenom	through,
krigets	the war's,war,
sjunde	seventh,
musikens	music,the music's,
berättat	told,
klubbarna	clubs,the clubs,
berättar	tells,
berättas	(as) told,is told,told,
korn	korn,barley,grains,
rester	residue,remains,residues,
dras	draw,preferred,make (assumptions, references),
drar	drag,earn,
inkomstkälla	income cold,source of income,was added to cold,
william	william,
drag	trait; characteristic; feature,move,characteristic,
mästare	master,champion,
matematiska	mathematical,
resten	the rest,rest,
jagar	hunts,hunting,
kors	cross,
närmaste	nearest,closest,
samarbetade	collaborated,collaboration,
enade	united,
medför	result,entails,means,
dvd	dvd,
officerare	officers,officer,
tunga	heavy,tongue,
heath	heath,
tillfälliga	temporary,
folkliga	popular,folk,
tungt	heavy,
svt	svt,
dvs	(det vill säga) namely that,d.v.s.,i.e.,
skyskrapor	high rise buildings; sky scrapers,skyscrapers,
stones	stones,
bonniers	bonnier's,bonniers,
höst	autumn,fall,
placera	position,place,
indiska	indian,
katt	cat,
företeelse	experience; phenomenon; feature,feature,phenomenon,
lutning	closing,angle,incline,
ge	to give,give,
tänker	thinking,
ga	ga,
go	go,
gm	by,
träd	into,tree,
kate	kate,
världsrekord	world record,
baron	baron,
uppgörelse	settlement,agreement,deal,
tillhör	belongs,belonging to,
flitigt	actively,frequent,
dröjde	slow,was not until,not until,
tänkandet	thinking,the way of thinking,
skildras	is depicted,depicted,
wave	wave,
rinner	running,flow,flows,
kommunismen	communism,
försvarsminister	minister of defence,
michael	michael,
ryan	ryan,
utbredning	distribution,distrubution,
tidszoner	time zones,
jönköping	jönköping,jonkoping,
stift	pin,diocese,
akut	urgent,acute,
oklart	clear,
socialdemokratiska	socialists,social democratic,
zh	zh,
derivator	derivative,derivatives,
mussolinis	mussolini's,mussolini,
honan	the female,female,
geologiska	geological,
visserligen	certainly,although,
början	top,beginning,
intervjuer	interviews,
singapores	singapores,singapore's,
kombination	combination,
kolonialism	colonialism,
geologiskt	geologically,geological,
svagare	weaker,weak,
kinas	china's,kinase,chinas,
erövringar	conquests,
hansson	hansson,
bjöd	offered,invited,
polen	poland,pole,
byttes	changed,was exchanged,
genombrott	breakthrough,
cell	cell,
experiment	experiment,
förhistoria	prehistory,
valen	the elections,elections,
gasen	gas,
utrikespolitiken	foreign policy,the foreign policy,
invigdes	inaugurated,
bindande	binding,
offentlig	public,published,
innerstaden	inner city,
händelsen	the occurence,event,
gåva	gift,
eminem	eminem,
vreeswijk	vreeswijk,
uppgick	total,was,
ryska	russian,
händelser	handelsar,happenings,events,
innebandy	floorball,
svenskans	the swedish language,swedish language,
västerut	west,westwards,westward; west,
chans	chances,chance,chanse,
överlevnad	survival,
tills	until the,until,
dopamin	dopamine,
uppfinningar	inventions,
arthur	arthur,
färöarna	faroe islands,the faroe islands,
vuxen	adult,
italienska	italian,
genetiska	genetic,
personen	person,the person,
utdöda	extinct,
genetiskt	genetically,genetic,
coldplay	coldplay,
kunde	could,
stärka	enhance,strengthen; bolster,
personer	person,persons,people,
jonathan	jonathan,
sjunger	sings,singing,
starten	the start,start,
mexikanska	mexican,
about	about,
invigningen	inauguration,the opening,
huxley	huxley,
misslyckades	failed,
släppte	released,
debutalbum	debut album,
släppts	released,
mottagaren	the receiver,the recipient,receiver,
guds	god,god's,
kenny	kenny,
utomstående	outside people; outsiders,outside,outsider,
linköpings	linkopingas,linköpings,linköping's,
halloween	halloween,
beslöt	resolved,decided,
studioalbum	studio album,
talat	spoken,spoke,
fördelningen	distribution,
talas	spoken,is spoken,
talar	speaks,talk,speak,
romantikens	the romanticism,romantick,romanticism,
tåget	train,the train,
kretsar	circuits,circles,circuitry,
tågen	train,the trains,
sovjetunionen	the soviet union,soviet union,
fälttåg	crusade,campaign,
ferdinand	ferdinand,
folkmängd	population size,population,
kronprinsen	crown prince,the crown prince,
oroligheter	unrest,
fara	danger,
uttalet	the pronounciation,pronunciation,
svenskar	swedish,swedes,
dödlig	lethal,mortal,
sena	late,
fars	father's,father,
utfördes	carried out,was carried out,preformed,
ringde	called,
österrikiska	austrian,
säljer	sells,
reagerar	react,reacts,
tillhöra	belong to,belonging to,
absint	absinthe,
artisterna	aristerna,artists,
encyclopedia	encyclopedia,
rörde	had something to do with,touched,was about,
kungliga	royal,
socken	parish,
högtider	holiday,feasts,
timmar	hours,
presidenter	presidents,president,
offentliga	public,
förstördes	destroyed,was destroyed,
någonting	nothing,anything,
fortsättning	continuation,continued,
presidenten	president,the president,
offentligt	public,publicly,
öarna	the islands,islands,
verklighet	true,reality,
belopp	amounts,amount,sum,
tränger	forces forward,cut in,penetration,
begick	commited,committed,
kyrkor	churche,churches,
insekter	insects,
allting	everything,
filosofiska	philosophical,
naturgas	natural gas,
konserten	the concert,concert,
zagreb	capital of croatia,zagreb,
ägna	baiting,spend,devote,
läror	teachings,
front	front,
konserter	conserts,concerts,
dikt	poem,
intäkterna	the revenues,proceeds,the revenue,
miniatyr|px|den	miniature,
hunden	the dog,dog,
kläder	clades,clothes,
university	university,
räckte	enough,handed,
finnas	found,(be) found,exists,
mode	fashion,mode,
förmågor	abilites,capacities,abilities,
modo	modo,
täcker	attacks,covers,
stadsparken	city park,stadsparken,city ​​park,
föreslogs	suggested,was suggested,proposed,
illuminati	illuminati,
globe	globe,
skolgång	school attendance,schooling,
 procent	percent,per,
stiger	rises,rising,
osmanerna	ottoman turks,ottomans,
apartheid	apartheid,
skov	forestry,episode,relapse,
skor	shoe,shoes,
special	special,
flyr	flees,escapes,
entertainment	entertainment,
förutom	besides; in addition to; aside from,except,
islamisk	islamic,
samarbetar	cooperate,cooperates,collaborates,
samarbetat	collaborated,collobrated,
max	max,
solsystem	solar system,
vinter	winter,
omfatta	cover,
torres	torres,
frånträde	relinquishment,withdrawal,
bilder	images,pictures,
lycka	happiness,good luck,
lida	sheath,suffer,
bilden	image,the image,
förstod	understood,
förbund	union,federal,league; alliance; union; compact; covenant,
kommunala	local,municipal,
livsmedel	food,
banor	paths,line,
times	times,
åter	again,undertake,
benämnas	named,entitle,entitled,
strida	conflict,fight,
tillgången	access,
tigrar	tigers,
austin	austin,
partierna	portions,political parties,
riksdagsvalet	parliamentary election,election to parliament,parliamentary elections,
ursprungsbefolkningen	the native population,indigenous people,indigenous population,
brandenburg	brandenburg,
centrum	center,
bedöma	judge; decide,assessment,
kategorihedersdoktorer	category of honorary degrees,
spaniens	spain's,
ipredlagen	ipred act,
attack	attack,
boken	paper,the book,
mao	mao,
dygnet	day,
infaller	no cells,falls,
final	final,finite, final,
zeeland	zealand,zeeland,
nilsson	nilsson,
belgiska	belgian,
hasch	hashish,
emellertid	however,
styrelseskick	form of government,government,
lista	list,
definierat	defined,
ben	bone,
definieras	defined,is defined,defines,
definierar	defining,defines,
arbetade	worked,
inbördes	relative,intermutual,
israelisk	israeli,
ber	ask,asks,
bet	bit,
julian	julian,
kvinnans	female,
hjärna	brain,
need	need,
bordet	the table,desktop,
varade	duration,lasted,
förra	last,former,
tredjedelar	thirds,
visor	songs,
förlorades	lost,was lost,
släkt	pettigree,family,
attackerna	attacks,the attacks,attack,
runorna	the runes,runes,
röst	voice,
förblev	remained,
jorge	jorge,
galleri	gallery,
regn	rain,
montana	montana,
genomslag	impact,breakthrough,
regi	direction,
tyskar	germans,
sändas	broadcast,be transmitted,sent,
nå	access,reach,
planerar	is planning,plan,planned,
skogar	forests,
långtgående	far-reaching,
platon	platon,platonic,
parker	parker,parks,
fiktiv	fictive,fictitious,
tolkien	tolkien,
fynden	finds; findings,findings,
försvara	research be,defend,defending,
skedde	was,
passa	take the opportunity,match,fit,
parken	park,the park,
hade	was,had,
basen	became,the base,base,
radioaktivt	radioactive,
baser	bases,
gemensam	joint,common,
härskare	ruler,
förbli	remain,
varit	has been,been,
partnern	partner,the partner,
aspekt	aspect,
psykologin	the psyhology,psychology,
boris	boris,
klassiska	classic,
inbördeskrig	civil war,
omloppsbana	orbit,
michigan	michigan,
förbjöd	forbade,forbid,
området	the area,area,
inflytelserika	influential,
klassiskt	classical,classic,
häst	horse,equine,
områden	areas,area,
unionen	union,the union,european union,
karriären	career,the career,
älskade	loved,loved; beloved,
gray	gray,
evolution	evolution,
processer	processes,
tillgång	access,
mohammed	mohammed,
grav	tomb,grave,
gran	spruce,
influensa	flue,influenza,flu,
också	also,
grad	grade,rate,
kvadratkilometer	square kilometer,square kilometers,
processen	process,the process,
vänt	turned,
sydafrika	south africa,
lätta	light,lighten,
västindien	caribbean,west india,
förband	units; formations; bound (themselves),bond,
neutralt	neutral,
korea	koreans,korea,
stats	state's,state,
tenn	tin,
lissabon	lissabon,lisbon,
flicka	girl,
gotiska	gothic,
staty	statue,
state	state,
företagets	the company's,the corporation's,
ken	ken,bank,
högra	right,
ersätta	replacing,replace,
sovjetiska	soviet,sovjet,
satsa	bet,
benämningen	the designation,the name,label,
merry	merry,
jobba	work,
befälet	the command,command,
distribution	distribution,
hits	hits,
innanför	inside,within,
synvinkel	angle,perspective,
vulkaner	volcanos,volcanoes,
framgångsrika	successful,successes,succesful,
trädde	met,entered,come into effect,
varierade	varied,
älskar	loves,
stratton	stratton,
framgångsrikt	successful,successfully,
partiklar	particles,
jersey	jersey,
uppsättning	equipment,set,
fördelar	advantages,share,advantage,
helsingfors	helsingfors,helsinki,
jim	jim,
opposition	opposition,
dominerande	dominating,dominant,
kategoribrittiska	category: british,category uk,
knst	knst,
leipzig	leipzig,liepzig,
johans	johan's,johan,
revolutionen	the revolution,revolution,
johann	johann,john,
kings	kings,king's,
sammanhang	connection,context,
christer	chris,christer,
willy	willy,
trycket	pressure,
sara	sara,
fokusera	focus,
äldre	old,older,
poet	poet,
påminde	reminded,
poes	poe,poe's,poes,
kingston	kingston,
vinci	vinci,
övertalade	over spoke,persuaded,
affärer	business,
spanska	spanish,
spaniel	spaniel,
spanien	spain,
humör	temper,mood,
strömningar	sentiments,tendencies,
kanarieöarna	canary islands,the canary islands,
 meter	metre,meters,meter,
erbjuda	offer,
reaktionerna	the reactions,reactions,
könsorganen	sex organs,the genitals,the reproductive organs,
utgjorde	made up,was,comprised; consisted of,
platons	platon's,plato,platos,
reaktion	reaction,reaction reaction,
vilkas	whose,
rysslands	russia's,
enkel	simple,plain,
feber	fever,
demo	demo,removed,
rättigheter	rights,
mysterium	mystery,
nordirland	north ireland,northern,
måleri	painting,
kategorikrigsåret	category war years,
alfabetisk	alphabetical,
revir	turf,territory,
reformationen	reformation,the reformation,
parti	party,batch,
instabil	unstable,
campus	campus,
varmed	whereby,
begav	went,went (to),traveled,
griffon	griffon,
dickens	dicken's,dickens,
korrekta	correct,
växjö	växjö,
flygbolag	airline,carriers,
anka	anka,duck,
nationens	the nation's,nation,
rankas	ranks,rank,
särskild	specific,particular,
införa	introducing,introduce,
eklund	eklund,
nämligen	namely,
spred	spread,
alperna	alps,the alps,
lagring	storage,
flickan	girl,the girl,
strömmen	current,the stream,
grenar	branches,
i	of,in,
kärleken	love,the love,
theodor	theodor,
europarådet	council of europe,european council,
onda	evil,
öga	eye,
störta	rush,crash,interfere,
sänds	sends,sands,sent,
sofia	sofia,
omkom	perished,died; was killed,died,
himmler	himmler,
förekommer	occurs,preferred is,
sända	transmitting,broadcast,send,
sände	sent,
vida	broad,wide,
jeff	jeff,
reducera	reduce,
natt	night,
nato	nato,
sweet	söt,
titta	see,watch,look,
bebyggelsen	building,human settlement,settlement,
jesper	jesper,
katolska	catholic,
utan	without,
sanning	true,truth,
vanligare	more common,
historia	history,
definitivt	permanent,unavoidable,definitely,
historik	history,
klassificering	classification,
loss	unstuck,off,
lincoln	lincoln,
lost	lost,
norges	norway's,
fernando	fernando,
martin	martin,
page	page,
regeringar	rings,governments,
lager	layer,
kolonierna	colonies,
vardagliga	ordinary,everyday,
pojkarna	boys,the boys,
library	library,
förlusterna	the losses,loss,
vardagligt	everyday,
förenklat	simplified,made easier,
omöjligt	impossible,
skorpan	crust,
peter	peter,
lagen	the law,law,
moskva	moscow,
skrifter	writings,
 km²	kilometres,
jugoslaviska	yugoslav,jugoslavian,yugoslavian,
hyser	has,accomodates,holds,
folkets	the people's,people,
slott	castle,
alliansen	the alliance,alliance,
fanns	was,
förde	led,out,
skriften	no.,writings,
broar	bridges,
hinder	obstacle,barrier,
motsättningar	contradictions,oppositions,frictions; clashes,
meddelade	informed; announced,announced,stated,
samlades	collected,gathered,were united,
journal	journal,jurnal,
reza	reza,
kromosomer	chromosomes,
halvön	peninsula,the peninsula,
småland	smaland,småland,
usas	usa:s,u.s.,
keramik	ceramic,ceramics,
freedom	freedom,frihet,
beslutade	resolved,decided,
samlats	collected,gathered; collected,
skrev	said,
polisens	police,the police's,
troligen	probably,likely,
synsätt	effects,viewpoint,
hävdade	argued,claimed,
mytologi	mythology,
betydelsefulla	significant,
glenn	glenn,
underjordiska	underground,
räddade	saved,
tendenser	tendencies,
längsta	maximum,longest,
utility	utility,
hammarby	hammarby,
pc	pc,personal computer,
museum	museum,
djävulen	devil,the devil,
realiteten	de facto,reality,
afrika	africa,
oändligt	infinity,infinitely,
heydrich	heydrich,
cricket	cricket,
north	north,
står	standing,star,stand,
instiftade	established,instituted,created,
neutral	neutral,
hn	hn,
ho	ho,
behov	necessary,
hc	h.c.,h.c,
ha	be,have,
he	he,
överens	in agreement,agree,
avled	deceased,died,
svarta	black,
stål	steel,
fysik	physics,
allierad	allied,ally,
dator	computer,
pippin	pippin pippin pippin,pippin,
komiker	comic,comedian,
förslaget	proposition,the suggestion,research team,
hästar	horses,
invandring	immigration,
bitar	bit,pieces,
farlig	dangerous,hazardous,
pelle	pellet,pelle,
ordbok	glossary,dictionary,
ibland	sometimes,
erik	erik,
själ	shawl,soul,
motsvarar	comparable,corresponds to the,corresponds,
eric	eric,
diego	diego,
omväxlande	varied,
sänktes	sunk,reduced,
moderaterna	the moderate,the moderates,moderates,
speciell	specific,special,
mineraler	minerals,
serveras	served,is served,
vulkaniska	vulcanic,volcanic,
canada	canada,
stat	state,
hittade	found,
liter	liters,
pontus	pontus,
revolutionära	revolutionary,
musikvideor	music videos,
stad	city,
musikvideon	music video,
resulterade	resulted,
stan	town,
bly	led,lead,
hjärnan	brain,the brain,
stam	strain,tribe,
etiken	the ethic,ethics,
förekomma	occur,be found,
inser	recognize,realizes,
klass	grade; class,class,
alkohol	alcohol,
simpson	simpson,
konsumtion	consumption,
hinner	reach it (in time),have time to,time,
felaktig	incorrect,false,error,
auktoritära	authoritarian,
protest	protest,
andra	second,other,
fredrik	fredrik,
flest	most,the most,
buddy	buddy,
likaså	also,as well,
upplagan	edition,
swan	swan,
kommersiellt	commercial,
kulturell	cultural,
bli	be,become,
kommersiella	commercial,
köpmän	traders,merchants,
gjordes	made,was,was made,
hemmet	home,the home,
kristendom	christianity,
östersjön	baltic,balticsea,
vasa	vasa,
åstadkomma	provide,create,achieve,
upplysningen	the enlightenment,enlightenment,
kända	known,
kände	felt,
examen	exam,degree,
disneys	disneys,disney,disney's,
behövdes	required,
försöka	try,attempt,
chokladen	the chocolate,chocolate,
avståndet	distance,the distance,
sydväst	southwest,
slogs	fought,was,
sexton	sixteen,
dagens	current,todays,
upp	up,
rollfigurer	roll model,role figure,characters,
force	force,
berlins	berlin's,berlin,
förstaplatsen	first place,
bröstet	chest; breast,breast,
dennes	his,
avfall	waste,
neo	neo,
nej	no,
kommissionen	commission,the commission,
unescos	unesco,
ned	down,bottom,
trodde	thought,
uppdelningen	partitioning; sectionalization; division; split (-ting),splitting,division,
new	new,
tätort	urban,conurbation,
ner	bottom,
ort	neighborhood,place,location,
med	with,
genomföra	perform,out,
men	but,
drev	pursued,drove,led,
vinden	the wind,wind,
pedro	pedro,
mer	more,
luther	luther,
geografiskt	geographically,geographic,
därpå	then,thereon,darpa,
oro	anxiety,worry,concern,
åka	go,
fyllde	completed,filled,
dubbla	double,
guide	guide,
kolonier	colonies,
geografiska	geographical,spatial,
dra	pulling,pull; (with)draw,
california	california,
magnusson	magnusson,
reste	stood,travelled,moved,
högtid	festival,festival; holiday,
£m	million pounds,
efterföljare	following,follower,successors,
rosenberg	rosenberg,
reagan	reagan,
atlanten	atlantic,the atlantic ocean,
inleddes	started,began,initiated,
fördelning	distribution,
soldat	soldier,
moral	morality,
berättelserna	the stories,stories,tales; stories,
prokaryoter	prokaryote,
gävle	gävle,
lennart	lennart,
provisoriska	provisional,
rockband	rock band,
bytet	the exchange,change,
oscar	oscar,
ljus	light,
nervsystemet	nervous system,the nervous system,
berlin	berlin,
upplevde	experienced,felt,
wikipedias	wikipedia,wikipedias,
ljud	sounds,noise,
köln	cologne,köln,
kategorikvinnor	category women,
flora	flora,
trots	although,despite,
procent	percent,per,
besittningar	holdings,possessions,
kapitalistiska	capitalistic,capitalist,
sundsvall	sundsvall,
kanadas	canada's,
erövringen	conquest,
tidskriften	the magazine,magazine,
abstrakta	abstract,
världskrigets	the world war's,world war,
förväntade	expected,
talets	the speechs,it means "decade" but would translate as "1950s", adding an s to the year.,century,
klitoris	clitoris,
konstitutionen	constitution,
tusen	thousands,
tidskrifter	magazines,periodicals,
risk	risk,
vänster	left,
satt	saat,sat,
nobelstiftelsen	nobel foundation,
bonaparte	bonaparte,
avrättningen	execution,the execution,
trött	tired,
begrepp	term,concept,
polis	police,
autonoma	autonomous,autonomic,
stilla	still,stationary,
tycktes	seemed,
orsakar	causes,
orsakas	caused,causes,caused by,
orsakat	caused,
utomeuropeiska	overseas,non-european,
gård	farm,house,
könsorgan	was organ,sex organ,genitals,
klarar	do,handle,
president	president,
orsakad	caused,induced,
indelat	divided,split,
medföra	bring,lead; result in, imply; entail,result,
indelas	divided,categorized,
indelad	divided,
medfört	resulted,led to,
låtskrivare	songwriter,song writers,
självklart	course,
indisk	indian,
ändra	change,
kvicksilver	mercury,quicksilver,witty zeal,
förfäder	ancestors,
fifa	fifa,
föreställningen	the idea,the concept,show,
panthera	panthera,
ibrahimović	ibrahimovic,
munnen	the mouth,mouth,
murray	murray,
föreställningar	performances,notions,
helena	helena,
buddhister	budhists,buddhists,
ovanstående	above,
listor	lists,
personal	personal,employed,staff,
förödande	devastating,
amerikanen	american,the american,
amerikaner	american,americans,
irans	iran's,
federationen	federation,the federation,
förstnämnda	first-named,aforementioned,first named,
förlängning	overtime; extension; prolongation,extension,
infektioner	infections,infection,
aston	överraska, undra,aston,
startat	started,
medlemmar	members,
downs	down,
stimulerar	stimulates,stimulating,
omgivning	surroundings,ambient,surrounding,
isen	the ice,
myntades	coined,was coined,
huvudrollen	the main role,leading part,
inledde	started,launched,
tillvaron	existence,life,the subsistence,
sida	website,page,side,
överraskande	surprisingly,
skeppet	the ship,nave,
side	side,
kammaren	chamber,the chamber,
bond	bond,
liga	compatible,league,
päls	fur,
mediet	medium,the medium,
medier	media,medias,
milan	milan,
aids	aids,
håret	hair,the hair,
kiev	kiev,
uppsala	uppsala,
årsåldern	age group,years old,
hänvisa	reference,refer,
talet	rate,century,
ihop	up,together,
talen	rate,years,
sluta	end,stop,
återfanns	was rediscovered,found,can be found,
venezuela	venezuela,
bestod	was,
foto	photo,
neutroner	neutrons,neutron,
larssons	larsson's,
normer	norms,standards,
stöds	supported,stood,is supported,
nietzsche	nietzsche,
nomineringar	nominations,
uppförande	code,construction,behavior,
folkvalda	elected,popularly elected,
faktum	fact,
iso	iso,
reinfeldt	reinfeld,reinfeldt,
representant	representative,
sökte	searched,
starta	start,startup,launch,
stewart	stewart,
gå	go,
nätet	net,the internet,
jordanien	jordan,
arrangeras	(is) arranged,arranged,arrange,
skalvet	quake,
leddes	passed,was led,
massiv	massive,
objektet	the object,object,
föreslagit	suggested,proposed,
girls	girls,
vikingatiden	vikings,the viking age,
förbi	past,past the,pass,
objekten	items,objects,the objects,
hollywood	hollywood,
någonstans	somewhere,nowhere,
representerade	represented,represent,
alfred	alfred,
åskådare	spectators,audience; viewer,
medeltiden	middle ages,
besegrades	defeated,
skaffade	acquired,aquired,took,
sabbath	sabbath,
grönwall	grönwall,gronwall,
symptom	symptoms,symptom,
hundar	dogs,
chef	head,
formell	formal,
kontrast	contrast,
antarktis	antarctica,antarctic,
street	street,
regissören	director,
härkomst	origin,provenance,
parter	party,sides,
troligtvis	probably,
bobo	bobo,
palace	palace,
stadsdelen	the district,district,
låta	let,
mina	my,mine,
modern	modern,
självständiga	independent,sjalvstandiga,
självständigt	independent,independently,independant,
triangel	triangle,
tecken	sign,characters,signs,
lämnar	leaves,
lämnas	left,
lämnat	left,
skildringar	scenes,description,descriptions,
tidiga	early,
monetära	monetary,
österrike	austria,
muskler	muscles,
förefaller	appear,it seems,appears,
tidigt	early,at an early stage,
tål	is resistant to,stand,can take,
blue	blue,
dessa	this,these,
bildar	serves as,form,
bildas	formed; made up (of),formed,
tåg	rail,trains,
bildat	formed,
mario	mario,
dödsfall	death,deaths,
luthers	luthers,luther's,luther,
vidsträckta	broad,wide; broad,
marie	marie,
typ	kind of,type,
diskuterats	been discussed,discussed,
maria	maria,
don	don,
utrustning	equipment,gear,
materiella	material,
talanger	talents,
dog	died,
slipknot	slipknot,
läsare	readers,reader,
points	point,
innersta	innermost,inner,
dos	dosage,
dop	baptismal,baptism,
kristen	christian,
långvariga	long,long-standing,
koppla	coupling,connect,
införde	enforced,introduced,
hjälper	helps,shows,
västeuropa	western europe,west europe,
befälhavare	commander,
liza	liza,
droger	drugs,
skyldig	responsible,guilty,
långvarigt	long-running,prolonged,long-standing,
nevada	nevada,
odling	cultivation,
krönika	chronicle,
anländer	arrive,arrives,
folkrepubliken	people's republic,people"s republic,
folke	folke,
helhet	entirety,whole,
monica	monica,
stycke	piece,piece; part; section,
meningar	sentences,
kollapsade	collapsed,
stop	stop,
stor	big; great,large,great,
stol	chair,seat,
strategiska	strategical,strategic,
präster	priests,
christopher	christopher,
stod	stood,
mönster	marks,
sandy	sandy,
earl	earl,
bar	bar,
bas	base,
existerar	exists,
skrivas	written,printed,
romerskkatolska	roman catholic,
existerat	existed,
anlades	founded,were built,was built,
bad	bath,
fokus	focus,
förändra	change; alter; replace,change,
gärningar	deeds,
anknytning	tie,link,related,
avvikande	different,deviant; divergent; different,
zonen	the zone,zone,
zoner	zones,
gunnar	gunnar,
vända	turn,habituated,
dittills	thus far,so far,
vände	reversed,turned,
turnén	turn,tour,tournament,
öppnade	opened,opening,
inledningsvis	initially,in the beginning,by way of introduction,
skrevs	written,was,
naturligtvis	course,off course,naturally,
skrift	no.,book,writing,
underart	subspecies,
sorts	variety,
göta	göta,
omkringliggande	surrounding,neighbouring,
smguld	swedish championship gold,sm gold,gold medal in the swedish championships,
artikel	article,
armeniska	armenian,
ondska	evil,
nationalister	nationalists,
bidragande	contributors,
kämpa	fight,
motto	motto,
regelbundet	regularly,regularily,
isotoper	isotopes,
fns	un's,tris,
regering	the government,government,
näringslivet	business,industrial life,economic life,
fördraget	the treaty,treaty,
fördragen	treaties,the compacts,
kol	charcoal,coal; charcoal,
ung	young,
ernst	ernst,
regelbunden	regular,
upptäcker	discoveries,discover,discovers,
atombomberna	atom bombs,the nuclear bombs,atomic bomb,
mellanrum	space,gap,
nationalförsamlingen	national assembly,
synsättet	approach,view,
avsikt	intention,intends,
interna	internal,
omstritt	controversial,
varmt	hot,warm,
erövrade	conquered,
studerat	studied,
blodkroppar	blood cells,corpuscle,
cyrus	cyrus,
varma	hot,warm,
tina	defrost,thaw,tina,
tillämpa	administer,implement,applying,
idol	idol,
minoriteten	minority,
betydelsefull	meningful,significant,
knutsson	knutsson,
igång	start,start up,
provinsen	province,the province,
utseende	appearance,
sällskapshundar	pet dogs,companion dog,
namnen	the names,names,name,
mindre	smaller,less,
etniskt	ethnical,ethnic,
azerbajdzjan	azerbaijan,azerbaijani,
blåvitt	blåvitt,bluewhite,blue and white,
etniska	ethnic,
pornografi	pornography,
paradiset	the paradise,paradise,
ix	4,the ninth,
förgäves	in vain,
albaner	albanians,
mexico	mexico,
kvinnor	female,women,
ip	ip,
sushi	sushi,
iu	iu,
it	it,
ii	(ii),
hämnd	revenge,
cant	cant,
djur	animals,animal,
im	im,
il	il,
in	in the context: recorded = spela (in),in,
colosseum	colosseum,
turner	tournament,
stoppa	stop,
konkurrensen	the competition,competitive,
vänstern	the left wing,left party,western,
make	make,husband,
producerats	produced,produced (by),
bella	bella,
västberlin	west berlin,
kommunistpartiets	communist party,the communist partys,the communist party,
roland	roland,
därmed	consequently,thus,therefore,
industriell	industrial,
makt	power,
benämningar	terms,names,
anglosaxiska	anglo-saxon,
atmosfären	atmosphere,the atmosphere,
försvarets	defense,forsvarets,the defence's,
dillinger	dillinger,
övriga	other,others,
kim	kim,
nicklas	niclas,nicklas,
folkrikaste	populous,people rich,most populus,
akademiska	academical,academic,
protesterna	protests,the protests,
nedan	below,hereinafter referred to as,
vetenskaplig	learn scientific,scientific,
sydamerika	south america,
glädje	joy,
dåvarande	then,formerly,
värmland	wermlandia,värmland,
roma	roma,
viktiga	important,
grannländer	neighbors,neighboring countries,neighboring lander,
facto	facto,
just	right,currently,just,
diameter	diameter,
jämför	compare,
sporting	sporting,
universitet	university,
psykos	phychosis,psychosis,
bollen	the ball,ball,
västeuropeiska	western european,
zon	zone,
human	human,
anders	anders,
beskriver	describes,
premiärminister	prime minister,
fysiker	physicist,physicists,
hävdar	states,assert,maintain,
bokstäver	letters,
troligt	likely,
hävdat	argued,claimed,
självstyrande	self-governing,independent,self-governance,
strax	soon,just,
royal	royal,
julen	julien,christmas,
memoarer	memoirs,
jules	jules,
friedrich	friedrich,
amerikas	america,america's,
harald	harald,
borgen	castle,bail,the castle,
komintern	komintern,comintern,
språkets	the language's,language,
arkitekturen	the architecture,architecture,
gustav	gustav,
behövde	did,needed,
rättegång	trial,steering wheel gang,
särdrag	special features,feature,features,
följaktligen	consequently,
utrikesminister	minister of foreign affairs,foreign minister,
tittar	looking; viewing; viewer,viewing,
författningen	constitution,
bekräftar	confirmed,confirms,
gustaf	gustaf,
trafikeras	served,trafficked,
trafikerar	traffic,frequent,
bekräftat	confirmed,
världsdel	continent,
sjöfarten	maritime transport,shipping,
medborgarskap	citizenship,
kommunerna	kommunera,municipalities,the municipalities,
släkting	relative,
intensiv	intensity,intense,
litauen	lithuania,
syrien	syria,
kemiska	chemical,
vattnet	water,the water,
kontinent	continent,
kunna	to,be able,
dead	dead,
befolkningen	the population,population,
uppmärksammades	attention,drew attention,
jupiter	jupiter,
befann	found,located,
kemiskt	chemically,
dominerade	dominated,
tappar	drop,lose,
statistik	statistics,
oralsex	oral sex,
hudfärg	color,
miljöproblem	environmental problem,environmental problems,enviormental problem,
teoretiska	theoretical,
hittades	was found,
däggdjuren	mammals,the mammals,
säsongerna	seasons,
shakespeare	shakespeare,
morden	murders,the murders,
värdefulla	valueable,valuable,value,
filmatiserats	cinematized,been filmed,screened,
benämns	designated,is mentioned,
knep	tricks,sleight of hand,
angrepp	attack,
burj	burj,
versioner	versions,
bolt	bolt,
härstamma	originate,stem,
burr	burr,
förkortas	shortened,abbreviated,reduced,
förkortat	shortened,abbreviated,
irländska	irish,
flyttat	moved,
fördelen	advantage,the advantage,
ljungström	ljungstrom,ljungström,
därutöver	in addition,addition,moreover,
maskiner	equipment,machines,
omröstning	vote,
mycket	very,much,
tillverkar	producing,makes,manufactures,
tillverkas	is made,manufacture,manufactured,
magazine	magazine,
ishockey	ice hockey,hockey,
strömmar	streams,flow,
grenen	the branch,branch,
förknippade	associated,
äktenskap	the marriage,marriage,
psykisk	psychic,mental,
romantiska	romantic,
français	francais,public,
grundades	founded,was founded,
jens	jens,
romulus	romulus,
orsak	reason,cause,factor,
down	down,
utbildning	education,eduction,education and training,
amsterdam	amsterdam,
havsnivån	sea level,
fastlandet	mainland,
estniska	estonian,
märks	notice,labeled,noted,
tennis	tennis,
könen	the sexes,equality,
bönder	farmers,
bolivia	bolivia,
märke	badge,label,
hyllade	celebrated,acclaimed,
form	form,
norrlands	northern sweden's,lapland's,norrland,
batman	batman,
ford	ford,
berg	mountain(-s),mountain,
civilisationer	civilizations,
japansk	japansk,japanese,
bero	depend,due,
bättre	better,
byggde	was,built,built, founded (on),
fort	fast,quickly,
tempel	temple,
spelade	played,
positiv	positive,
slaviska	slav,slavic,slavonic,
flickvän	girlfriend,
åriga	-year,year,
regeringen	the government,government,
båten	vessel,the boat,boat,
skelett	skeleton,
månens	the moon's,the moons,moon,
beteckningen	the label,designation.........,designation,
avsnitt	section,part,episode,
phil	phil,
petit	petit,
uttryckligen	explicitly,specifically,
handelspartner	trading partner,
tosh	tosh,
kanske	may,
primtal	prime number,
byggnaden	building,the building,
vista	vista,
handen	the hand,hand,
handel	commercial,trade,
kunnat	could,could have been,been,
svärd	sword,
betala	pay,
digital	digital,
betalt	charge,
marxism	marxism,
kungamakten	monarchy,the monarchy,
sades	said,was said,
överenskommelse	deal,arrangement,
frodo	frodo,
exporten	exports,the export,
jones	jones,
drivs	driven,run,powered,
accepterade	accepted,
engagemang	commitment,
riktad	directed,
ökande	increasing,rising,
fss	fss,
expandera	expand,
skuggan	shadow,the shadow,
riktas	directed (at),direct,target,
riktar	targets,target,
milt	mild,
armar	arms,
bomben	bomb,the bomb,
telefon	telephone,
tredje	third,
mild	mild,soft,
bomber	bombs,
vikingarna	the vikings,
marissa	marissa,
dä	the elder,with,
imperiet	the empire,empire,
avbrott	break,breaks,
uppdelning	division,partitioning,playback,
petersburg	petersburg,
dö	die,
lissabonfördraget	treaty of lisbon,lisbon treaty,
me	me,
illa	bad,
din	yours,your,
fackföreningar	unions,
dig	up,
trenden	trend,the trend,
afrikansk	african,
anna	anna,
dit	there,where,
spets	edge; top,tip,point,
bulgarien	bulgaria,
olympia	olympia,
ville	wanted (to),did,wanted,
malmö	malmö,malmo,
diskografi	discography,
villa	house,villa,
slagit	held,beaten,
reklamen	the commercial,commercial; ad; advertisment,advertising,
invandringen	immigration,
rymden	space,
utlösning	release,ejaculation,trigger,
hästen	the horse,
bakom	behind,
afghanistan	afghanisthan,afghanistan,
viktig	major,important,
kokain	cocaine,cocain,
föredrog	prefered,preferred,
bibliotek	library,
lönneberga	lönneberga,lonneberga,
somalia	somalia,
international	international,
madagaskar	madagascar,
avsluta	finish,exit,
nationalismen	nationalism,
tibet	tibet,
henry	henry,
högkvarter	headquarters,head quarter,
avsaknad	absence,
kommun	local,municipality,
beskrivits	described,
boy	boy,
diagnoser	diagnoses,
canadian	canadian,
institute	institute,
bor	lives,
främst	foremost; primarily; chiefly,all,primarily,
gyllene	golden,golden; gilded,
vietnamesiska	vietnamese,
bok	book,
mängder	amounts,amount,
extrem	extreme,
mänsklighetens	humanity's,humanities,
bolivianska	bolivian,
diagnosen	diagnosis,the diagnose,
departement	departement,department,
sporter	sports,
enorma	enormous,
utövar	exercises,carrying,exercise,
utövas	is practised,exerted,exercised,
världshälsoorganisationen	world health organization,
asiatiska	asiatic,asian,
sporten	the sport,sport,port,
religionsfrihet	freedom of religion,religious freedom,religion,
östasien	east asia,
platån	sycamore,the plateau,plateau,
skräck	fear,horror,
franco	franco,
hemmaarena	home ground,home field,
tennisspelare	tennis player,
socialister	socialists,
maya	maya,
peru	peru,
kristian	kristian,
statsmakten	the government,power,government,
left|px	left px,
österrikeungern	oster kingdom hungary,austria-hungary,
detaljer	details,
avsattes	deposited,dismissed,
brukade	used to,used,
ögon	eye (-s),eyes,
kemisk	chemical,
fartyget	vessel,ship; vessel,boat,
fly	escape,
hända	may,
hände	happened,
tokyo	tokyo,
mästarna	the champions,champions,the masters,
soul	soul,
träffades	met,was met,reached; met,
vittnen	witnesses,
akademien	the academy,academy,riksdagens,
präglade	characterized,
anslutna	affiliated,connected,
bristande	lack of,lack,wanting,
sökt	pending,searched,
ulf	ulf,
hiroshima	hiroshima,
crazy	crazy,
kenneth	kenneth,
uruguay	uruguay,
winston	winston,
agent	agent,
bemärkelse	meaning,sense,
skadades	damaged,was wounded,
beatles	beatles,
council	council,
dennis	dennis,
kunglig	royal,
pink	pink,piddle,
diskuterades	discussed,
oslo	oslo,
engelsmännen	english people,the english,the british,
varor	products,
ekonomiska	economic,economical,
till	to,
gitarrist	guitarist,
nya	new,
nye	new,
mat	food,
regeringstid	term of government,term of government; term of office,reign,
may	may,
överensstämmer	conform,agree,match,
uppföljare	sequel,
fotboll	football,
läkare	doctors,doctor,
maj	may,
upphört	ceased,left the association,end,
man	is,one,
asien	asia,
johnson	johnson,
kulturella	cultural,
sådana	such,
eng	eng.,
q	q,
tala	speaking,speak,
block	block,
basket	basketball,
romantiken	romance,romanticism,
undantag	exception,except,
sådant	such,
lsd	lsd,
bussar	bus,
bevisa	prove,
alfabetet	alphabet,the alphabet,
städerna	urban,the towns,
gällde	applied,applied to,was,
sällsynta	rare,
moralisk	moralic,moral,
huvudsak	in principal; chiefly,mainly,main thing,
lyrik	poetry,
motståndet	the resistance,the resistence,
verksam	active,effective,
landskap	province,landscapes,landscape,
juryn	the selection panel,the jury,jury,
sekter	sects,
inkomster	revenue,income,
äkta	genuine,married,authentic,
rasen	breed,the race,
policy	policy,
växte	grew,grow,
main	main,
texas	texas,
lägst	lowest,lowermost,
steget	step,
kräver	requires,
janeiro	janeiro,
domstolar	courts,
försörjning	sustention,sustentation,supply,
sibirien	siberia,
leds	led by,passed,
vindkraft	wind power,wind,
färg	colors,colour,
uppskattning	appreciation,estimated,
leda	lead,
villkoren	the terms,conditions,
rock	rock,
föremål	object,subject,
tysklands	germany's,germanys,
guevara	guevara,
latin	latin,
tacitus	tacitus,
hellre	rather,more preferably,
söner	sons,
vattendrag	water,streams,watercourse,
avkomma	progeny,offspring,
girl	girl,
dianno	di'anno,dianno,
saudiarabien	saudi arabia,
enastående	exceptional,outstanding,
jackson	mrs. jackson,jackson,
håkansson	hakansson,håkansson,
avrättningar	execution,executions,
pamela	pamela,
områdena	the areas,areas,
tronföljare	heir,heir apparent,successor,
kattdjur	felidae,cat,
valdes	representatives',selected,chosen; elected,
premiären	premiere,premier,
ansiktet	face,
monster	monster,monsters,
romani	romani,romany,roma,
konstnär	artist,
chiles	chiles,chile's,
tomt	empty,blank,
ajax	ajax,
snabbast	fastest,
brooke	brooke,
kognitiva	cognitive,
ord	word,words,
tunnelbanan	subway; tube; underground,the subway,metro,
keith	keith,
verkade	did,appeared to,were active, worked, was active,
gott	good,practically; good,
anledning	reason,
preventivmedel	contraceptives,
självmord	self-killing,suicide,
uppvisar	shows,
rankningar	ranking,rankings,
vision	vision,
stängdes	closed,
kraftig	strong,
egentligen	really,actual,actually,
first	first,
centrala	central,
grupperna	groups,
intryck	impression,appearance,
uttalanden	statements,
här	this; here,is,here,
rachel	rachel,
folklig	popular,folk,
biografen	the cinema,movie theater,cinema,
centralt	central,centrally,
skapandet	creation,the making,
kommunism	communism,
grundämnet	the element,element,
missnöje	dissatisfaction,
homogen	homogenous,
visar	is,shows,
består	consists of,beasts,exists,
västbanken	the west bank,westbank,
grundämnen	elements,
individ	individual,
örebro	Örebro,
öronen	lugs,the ears,
besluten	decisions,
anus	ass,anus,
köpenhamns	copenhagen,copenhagen's,
fysiska	natural,physical,
fysiskt	physically,physical,
danny	danny,
löstes	solved,dissolved,
drevs	concentrated,was driven,
beslutet	the decision,
konkreta	specific,concrete,
fiender	enemies,
fienden	enemy,the enemy,
medlemmarna	members,the members,
lugn	calm,
jordytan	earth's surface,earth crust,
fordon	vehicle/-s,vehicles,vehicle,
inträde	entry,
marklund	marklund,
jämlikhet	equality,
stadsdelar	districts,city districts,neighborhoods,
marijuana	marijuana,
större	greater,bigger,
formerna	forms,
tänder	teeth,
orsakerna	the causes,
kevin	kevin,
adeln	nobility,
nikola	nikola,
politiska	politic,political,
förälskad	in love,
menas	mean,means,
skulptur	sculpture,
centralbanken	centralbank,central bank,
potential	potential,
politiskt	political,
performance	performance,uppträdande,
centralstation	central station,
magnetiska	magnetic,
channel	channel,
norman	norman,
normal	normal,
hertig	duke,
dagbladet	daily paper,dagbladet,
fotografier	photographs,
halvan	the half,half,
politisk	political,
teoretiskt	theoretic,theoretical,
mordet	the murder,murder,
arbetat	worked,
queens	queen,
över	of,over,
visades	was,showed,
otaliga	countless; endless,countless,
lojalitet	loyality,loyalty,
drottning	queen,
grammatik	grammar,
österut	eastwards,east,
kontrolleras	is controlled,controlled,
kontrollerar	controlling,controls,controls; controlling,
ungdom	youth,
civilisationen	civilization,
show	show,
adolfs	adolf's,adolf,
uranus	uranus,
tidigast	the earliest,
or	or,
generalsekreterare	the secretary-general,secretary general,
samlingsalbum	compilation album,compilations,
helig	holy,
dick	dick,
historier	stories,history,
passande	fitting,suitable,matching,
historien	history,
black	black,
karolinska	karolinska (institute for medicine),caroline,
experimenterade	experimented,
ges	given,be given,
ger	gives; is giving,give,gives,
raser	races,species,
kulturellt	culture,cultural,culturally,
konsolen	bracket,
motsvarande	corresponding to,corresponding,
skådespelare	actor,
inspelningarna	recordings,
landets	the country's,its,
katla	katla,katla (fictive dragon in the classic "bröderna lejonhjärta"),
vintergatan	milky way,the milky way,
firade	celebrated,
ledaren	leader,conductor,
gen	gene,
beskyddare	protector,patron,
himmlers	himmlers,himmler,
mattis	mattis,
bengtsson	bengtsson,
statistiska	statistical,
tsaren	the czar,czar,the tsar,
spridda	spread,scattered,
europacupen	euro (-pean) cup,european cup,
miley	miley,
tolfte	twelth,twelfth,
relativt	relative,relatively,
sämre	poor,
sekulära	secular,
fokuserar	focuses,focus,
nazisterna	the nazis,nazis,
toppade	topped,
relativa	relative,
sean	seab,sean,
slöt	joined (in peace),closed,
utgiven	published,
menat	meant,
menar	mean,means,
kandidater	candidates,
försvarsmakten	national defense,national defence,armed forces,
döden	death,
vanns	was won,(was) won,
människan	the human,man,people,
söndagen	sunday,
personligt	personal,private,
världskriget	world war,
gaga	gaga,
människas	human's; man's,human,
personliga	personal,
förenta	united,
august	august,
 °c	celsius,
ju	the,the more,
tur	turn,tour,luck,
forskaren	researcher,
jr	jr.,junior,
åker	go,treats,field; going,
timme	hour,
tum	inch,inches,
fick	got,was,
signaler	signals,
lexikon	lexicon,
ja	yes,
ministrar	ministers,
rugby	american fotboll,rugby,
ån	on,from,the river,
utvalda	selected,selected; chosen,
tour	tour,
åt	to,for,
ås	ridge,site,
år	the year,year,
vätska	fluid,liquid,
naturresurser	natural resources,
jobb	job,work,
tryck	press,pressure,print,
vilja	will,like,
århundraden	centuries,
cancer	cancer,
statschefen	the head of state,head of state,
syntes	synthesis,
grundare	founder,
territorium	state,territory,
mätningar	measurements,measurments,
ryggen	the back,back,
barry	barry,
överföra	transmit,transfer,
bildats	formed,had formed,created,
kirsten	kirsten,kristen,
industrin	industry,
västliga	western,
utsatta	exposed,
mars	march,
överförs	is transferred,transfered,
plötsligt	suddenly,sudden,
marx	marx,
mary	mary,
kultur	culture,
flaggan	the flag,flag,
cobain	cobain,
partido	partido,
avskaffa	abolish,
bmi	bmi,
dvärghundar	miniature dogs,
spelfilmer	motion pictures,feature film,feature films,
klädsel	cover,
meningen	sense,
fortsatt	further,continued,
sound	sound,
metall	metal,
dragit	drawn,dragged,preferred,
uppstod	developed,was,
kategorimän	category: men,category men,
insåg	realized,
nionde	ninth,
sahara	sahara,
intressanta	interesting,of interest,
uppmanade	urged,encouraged,
liknande	similiar,similar,
sydkorea	south koreans,south korea,
hålls	maintained,maintaned,is held,
par	pair,
upplagor	editions,the edition,issues,
jesu	jesu,jesus,
edwin	edwin,
lava	lava,
hålla	hold,keep,
röka	smoking,smoke,
stött	met,supported,
pan	pan,
samt	also,as well as,
tidvis	times,
hösten	fall,the fall,the autumn,
running	running,
kuba	cubans,cuba,
teknisk	technical,
lösningar	solutions,
sömn	sleep,
markus	marcus,
fattas	taken,
bang	bang,
wahlgren	wahlgren,
identifiera	identification,
gates	gates,
münchen	munchen,munich,
bebyggelse	settlement,settlements,habitation,
privatliv	private,
reaktionen	reaction,the reaction,
dinosaurierna	dinosaurs,dinasaurs,
skapelse	creation,
väst	west,the west,
byggnad	building,
reaktioner	reactions,
våld	violence,force,
jakten	the hunt,hunt,
ideologiskt	ideologically,ideological,
grannländerna	neighbors,neighbouring countries,
bowie	bowie,
livstid	lifetime,life span,
programledare	host,
gotland	gotland,
ideologiska	ideological,
tros	belived,believed,
motverka	prevent,counteract,counter,
trä	wood,
möter	meets,meet,
vintern	the winter,winter,
schwarzenegger	schwarzenegger,
underarten	subspecies,sub species,
mån	concerned,mon,
mor	mother,
haft	had,
prägel	character,mark,
mot	against,
kategori	category,
jakt	hunt,hunting,
temperatur	temperature,
mon	mon,
underarter	sub-species,subspecies,
baltiska	baltic,
kollektiv	collective,public,
mod	courage,mod,
christina	christina,
adams	adams,
födda	born,
började	started,began,
födde	gave birth too,born,
jordbävningar	earthquakes,
manhattan	manhattan,
mänsklig	human,
sågs	observed,seen,was observed,
göran	göran,request,
bipolära	bipolar,
göras	made,be made,be made through,
rikskansler	chancellor,
kategorisveriges	category sweden,
joan	joan,
feodala	feudal,
konspirationsteorier	conspiracy theories,
förs	out,led,rapids,
jordbruket	agriculture,the agriculture,
lotta	raffle,lotta,
fört	led,lead,
sudan	sudan,the sudan,
reportrar	reporters,
föra	pre,lead,
före	ahead (of), before,present,before,
ända	as far as,up,
demokratisk	democratic,
traditionell	traditional,conventional,
ände	end,
moderata	moderate,moderates,
vistas	live,present,
förlust	loss,
londons	london's,
framstående	prominent,
olof	olof,
akon	akon,
tongivande	influential,
tillverka	producing,
sjätte	sixth,
celler	cells,
island	iceland,icelandic,
allians	alliance,
metaforer	metaphores,metaphors,metafor,
lands	land,on land,
lagarna	the laws,
retoriken	rhetoric,
auschwitz	auschwitz,
kort	short,
arvid	arvid,
wilde	wilde,
beskrivas	described,be described,
einstein	einstein,
mark	ground, soil, territory,ground,
intellektuella	intellectuals,intellectual,
floderna	floods,the rivers,rivers,
fullständigt	completely,full,
gravid	pregnant,
behandling	treatment,
varelse	creature,
emellanåt	once in a while,occasionally,
anfalla	attack,
välmående	healthy,well-being; affluent,prosperous,
fullständiga	full,complete,
kvinnlig	females,female,
tillfälligt	temporarly,temporary,
eget	own,
inletts	started,initiation,initiated,
utbredd	widespread,spread,
birger	birger,
härifrån	from here,here,
e	e,
egen	own,
tävlingen	competition,contest,
vhs	vhs,
exemplar	copies,example,
bibliografi	bibliography,
manuel	manuel,manual,
verkliga	real,fair,
identifierade	identified,
humanismen	humanism,
parlament	parliament,
håkan	håkan,chin,
följde	followed,
youtube	youtube,
manliga	male,
öns	the islands,island's,
prestigefyllda	prestigious,
skriven	written,
pompejus	pompey,pompejus,
arabiska	arabic,arabian,
goebbels	goebbels,geobbels,
film	film,
diktaturen	dictatorship,
again	again,
genrer	genres,
effekt	effect,power,
istanbul	istanbul,
spåren	the tracks,tracks,wake,
rubiks	rubiks,rubik's,
muren	wall,
produktiv	productive,productivity,
stannade	stayed,
spåret	groove,
genren	genre,
faktorer	factors,
däremot	on the contrary,however, on the contrary,however,
ordna	arranging,arrange,
profet	prophet,
ungarna	the kids,kids,the young,
förändrade	changed,
rykten	rumors,
ledning	conduit,guidance,
henriks	henry,
kyros	cyrus,
världsliga	worldly,
medicinska	medicinal,medical,
araberna	arabs,
palestinska	palestinian,
uppfostran	upbringing,
medicinskt	medical,
kuwait	kuwait,
snabbaste	rapid,fastest,
begå	commit,
resolution	resolution,
åtskilda	separated,segregated,separate,
mellanöstern	middle,the middle east,middle east,
vila	rest,
socialismen	the socialism,socialism,
inspirerat	inspired,
dollar	dollar,
vill	will,to,want,
hindrar	prevent,stop; prevent,prevents,
ingripande	negative,intervention,
inspirerad	inspired,
liam	liam,
levern	the liver,liver,
sund	healthy,narrow,sane,
symbolen	the symbol,
lugna	reassure,calm,
rwanda	rwanda,
symboler	symbols,
skydda	protect,protection,
skriver	write,type,
seriens	series,
kasta	discard,throw,
avhandling	treatise,thesis,
handlade	dealt with,was (about); traded,was,
israeliska	israeli,isrealic,
fall	where,
ramen	frame,
stödja	support,
ramel	ramel,
kulminerade	culminated,
ansvarig	charge,
miljoner	milions,one million,millions,
båtar	boats,
snuset	snuff,the snuff,
suttit	been,sat,
ockuperades	occupied,
cornelis	cornelis,
massor	lots,(in) masses,tons,
växthuseffekten	the greenhouse effect,greenhouse effect,
intressant	interestingly,of interest,
material	material,materials,
abc	abc (swedish news program),abc,
danmark	denmark,
publik	audience,public,
östtysklands	east germany's,osttysklands,
public	public,
lärare	teacher,
långhårig	rough,long haired,long-haired,
bebott	inhabit,inhabited,an inhabitated,
närhet	close,proximity,closeness,
vald	elected,selected,
jonas	jonas,
free	free,
benen	legs,
valt	chosen,selected,
sångare	singer,
historiker	historians,
jackie	jackie,
airport	airport,
uppslagsverk	encyklopedia,encyclopedia,
alexandria	alexandria,
ive	i've,
sjukhuset	the hospital,hospital,
africa	africa,
släktingar	relatives,
enat	united,
rösterna	votes,the votes,
författaren	the author,author,
hyllning	tribute,tribute; homage,
eye	eye,
torrt	dry,
utmärkelsen	award,the award,
innebar	meant,was; meant; entailed,was,
utmärkelser	commendations,awards,
torra	dry,
landet	state,the country,
diamond	diamond,
människa	human,man,
romersk	roman,
koma	coma,
brist	lack,non,failure; lack of,
tillkommer	reside,will be,will be added,
hundraser	breed of dogs,alternative strains,breeds,
skivor	plates,records,
berätta	tell,
vladimir	vladimir,
der	where,german word,
des	des,
det	is,it,dent,
roosevelt	roosevelt,
utsläpp	emission,emissions,
bron	bridge,the bridge,
del	part,
lindgren	lindgren,
den	it,
lagerlöf	lagerlof,lagerlöf,
befintliga	current,existing,
samtliga	all,
hastigt	rapidly,fast,
latinets	latin,the latin,the latin's,
sovjetunionens	soviet union's; soviet's,soviet union,
betoning	stress,
samhälle	society,
sjukdom	illness,disease,
medförde	resulted,brought,led,
födseln	birth,the birth,
sträng	string,strang,
robinson	robinson,
protein	protein,
makten	power,the power,
hämta	retrieve,fetch,
stil	type,
psykotiska	psychotic,
georgien	georgia,
stig	stig,path,
verkligheten	real,reality,
blad	leaves,leaf,
försvinner	disappears,disappearing,disappear,
primära	primary,
vikten	importance,weight,
makter	powers,
rastafari	rastafari,rastafarian,
avtalet	the treaty,the contract,agreement,
pettersson	pettersson,
laboratorium	laboratory,
ännu	even,still,yet,
judiska	jewish,
huvudkontor	central office,headquarters,
ligger	lies,is,
vatten	water,
rastafarianer	the rastafarian,rastafarian,rastafarians,
rockgrupper	rock groups,rock group,rock bands,
facebook	facebook,
beredd	ready (to),prepared,
konservatismen	conservatism,
civila	civil,
inåt	inwards,inwardly,
uppgav	said,
nordsjön	north sea,
officiella	official,
latinamerika	latin america,
fältet	the field,field,
förmågan	the ability,
göra	do,do; doing,
försäkra	insure,make sure,assure,
gradvis	gradually,progressively,
tvåa	second,
same	lapp,sami,
mörka	dark,
görs	is,made,is made to,
officiellt	official,officially,
människans	humans,mankinds,human,
längden	the length,length,lenght,
diskussion	discussion,
wilhelm	wilhelm,
edmund	edmund,
inbördeskriget	civil war; civil war,civil war,
epok	epoch,
odlade	grew,cultured,
saknades	lacked,missing,
trossamfund	religious community,faith community,religious communities,
suverän	terrific,supreme,sovereign,
good	good,
träffar	meets,hits,
ställas	set,be set,prepared,
planerna	the plans,plans,
fängelse	prison,
sexuellt	sexual,
oxford	oxford,
skrifterna	scriptures,
association	association,
toronto	toronto,
robbie	bobbie,robbie,
kungarna	the kings,kings,
namibia	namibia,
out	out,
byggt	building,built,
anslöt	joined,
trådlös	wireless,
house	house,
energy	energy,
hard	hard,
flytta	move,
öron	ear,ears,
förenade	united,
energi	energy,
perry	perry,
sanningen	truth,the truth,
östman	Östman,
oftast	usually,most often,
infrastrukturen	infrastructure,the infrastructure,
ölet	the beer,beer,
forskning	research,
perro	perro,
förföljelser	persecution,pursuits,persecutions,
fullständig	full,complete,n/a,
konflikt	conflict; strife,conflict,
prins	prince,
lawrence	lawrence,
strömning	flow,
eventuella	any,eventual,
blekinge	blekinge,
uralbergen	the ural mountains,urals,
eventuellt	eventually,possibly,
viken	gulf,
helsingör	helsingor,elsinore,helsingör,
inflationen	inflation,
investeringar	investments,
finland	finland,
jordens	earth,
utöver	addition,
fått	was given,with,
styre	governance,rule,
legenden	legend,
ensam	alone,
styra	controlling,steer,
top	top,
sjunkande	sinking; decreasing,decreasing,
dont	do,
säkerhetsråd	security,security council,
treenighetsläran	doctrine of the holy trinity,trinity,school of trinity,
snarast	rather,as soon as possible,
juridiska	juridical,legal,
carter	carter,
lidande	sufferer,
kom	came,
diskriminering	discrimination,
gator	streets,
kon	group,
åtta	eight,
observationer	observations,
förhindrar	prevents,prevent,
kategoriasiens	category of asia,
costa	costa,
kardinal	cardinal,
järnvägar	failways,rail,railways,
triangeln	triangle,the triangle,
part	party,
gudarna	the gods,
domstolen	court,the court,
direkta	direct,
matteusevangeliet	gospel of matthew,book of matthew,
följden	the result,the cause,result,
fattiga	poor,
knapp	scarce,button,bare,
proteinerna	the proteins,proteins,
ö	island,o,
personens	person,the persons,the person's,
börjar	starts,starts to,start,
hellström	hellström,hellstrom,
baháí	baha'i,bahá'í,
avtar	declines,avatar,
självständig	independent,independently,independant,
följder	impact,consequences,
följdes	followed,was followed,
rikedom	riches,wealth,
börjat	started,begun to,begun,
försökte	try,tried to,tried,
bränsle	fuel,
gjord	made,
flertalet	most,several,majority; plurality,
gjort	made,done,created,
mountain	mountain,
hundratals	hundreds of,hundreds,
mussolini	mussolini,mossolini,
infrastruktur	infrastructure,
caesar	caesar,
genast	at once,immediately,
taktik	tactics,tactic,strategy,
inkomsterna	the incomes,the income,revenue,
dramatiskt	dramatic,dramatically,
skjuta	delay,postpone; shoot,
militärt	military,militarily,
patterson	patterson,
krafter	forces,
gillade	liked,approved; liked,
niclas	niclas,
kraften	the force,power,
utbrott	outbreak,outbreaks,
samtidigt	while,simultaneous,
organiserade	organized,
högt	high,highly,
ko	co,cow,
km	km,kilometers,
kl	hr,at,o'clock,
kr	kronas,
liechtenstein	liechtenstein,
organisk	organic,
organism	organism,
thomas	thomas,
venedig	venice,venedig,
kvalitet	quality,
bergman	bergman,
relation	ratio,relation,
utveckla	develop,developing,
fina	beautiful,fine,
nämns	mentioned,
antagit	adopted,presumed,
konto	account,sign,
undre	lower,
wallenberg	wallenberg,
medverka	take part,participate,
världens	the world's,the world,the worlds,
tionde	tenth,
förbudet	ban,the union,
avseende	regard,for,
blomstrade	flourished,
typiskt	typically,typical,
nationalpark	national park,
kristina	kristina,
notation	notation,
beslutar	decides,
vänskap	friendship,
express	express,
beslutat	resolved,decided,
förklarat	explained,declare,
typiska	typical,
förklarar	explain,explains,
gamla	ancient,old,
husen	housing,the houses,
skickas	is sent,sent,any,
skickar	sends,send,
brukar	usually,used to,
wallander	wallander,
gamle	old,
uttrycket	the expression,expression,
uttrycker	express,expressing,express (-es),
flykt	escape,
huset	housing,the house,
svarar	responds,
somrar	summers,
stadium	stage,
styrdes	was guided,governed,ruled,
suveränitet	sovereignty,
rollfigur	character,
godkännas	approved,pass on,be approved,
höglandet	highlands,the highland,
tengil	tengil,
fann	found,
rovdjur	predator,predators,
fans	fans,
landsbygden	rural,rural area,
champagne	champagne,
romarriket	roman empire,the roman empire,
bildandet	setting-up,formation,establishment,
professionella	professional,
framförs	is presented,performed,
framfört	expressed,presented,
rörelserna	the movements,movement,
kritiserades	critisized,critizised,
framföra	express,convey,
skivorna	the records,records,plates,
medlem	member,
musklerna	muscles,the muscles,
statligt	state,governmental,
vuxit	grown,
praktiskt	convenient,
statliga	state,
restaurang	restaurang,restaurant,
baltimore	baltimore,
romska	romani,roma,
beta	graze,beta,
globala	global,
kroatiens	croatia's,croatias,croatian,
förklaring	explaination,explanation,statement,
point	point,
folkmord	genocide,
karaktären	the character,character,
andas	breath,breathes,
karaktärer	character,characters,
således	hence,thus,
tennessee	tennessee,
globalt	globally,global,
behöll	kept,retained,
försäljningen	sales,
lyfta	lift,
våningar	floors,storeys,
laos	laos,
bestämde	determined,chose,
inför	before,
bengt	bengt,
popularitet	popularity,
gav	gave,
effektiva	effective,
gas	gas,
vana	familiar,used,habit,
kalmar	kalmar,
effektivt	effective,
trupperna	troops,the troops,
detsamma	the same,same,
bild	picture,image,
motorväg	freeway,highway,
åtalades	was charged,was prosecuted,charged,
spridning	diffusion,distribution,proliferation,
bill	car,
döptes	renamed; named,renamed,baptised,
portugal	portugal,
arenan	arena,the arena,
elektronik	electronics,
påbörjade	started,
monroe	monroe - it's a persons name,monroe,
rederiet	the shipping company,the company,shipping company,
dödat	killed,
granska	examining,review,exam,
sjuk	ill,disease,
dödar	kill,kills,
dödas	put to death,killed,
hamna	end up,end,
motståndaren	the opponent,adversary,opponent,
administrationen	administration,
dödad	killed,
tyder	indicates,
sittande	fitting,appointed,sitting,
development	development,
övertogs	were taken,overtaken,
skotska	scotland,scottish,
syd	south,
konstnärliga	artistic,
syn	sight,view,
jerusalems	jerusalem's,
moment	step,
kallades	was called,called,summoned,
parentes	brackets,
avsett	avset,regard,intended,
nämnde	mentioned,said,
småningom	when the time comes,eventually,
tillbehör	sides,condiments,accessory,
nämnda	said,
kungariket	kingdom,the kingdom,
noll	zero,
kapitel	chapter,
albanien	albania,
jorderosion	earth erosion,soil erosion,
ministerrådet	minister counsellor,ministers,
värme	heat,thermal,
skott	bulkheads,round,shots,
albanska	albanian,
norrland	norrland,northern,
simmons	simmons,
bibeln	bible,
kommunister	communists,
juventus	juventus,
halvt	half,
organization	organization,
verkställande	executive,
passerar	passes,pass,
struktur	structure,
senaste	last,
billboard	billboard,
alternativt	alternatively,alternative,
sju	seven,
world	world,
analytiska	analytical,
alternativa	alternative,
tropisk	tropical,
sektion	section,
sparta	spartans,sparta,
administrativt	administrative,administratively,
monarkin	monarchy,the monarchy,
dömd	sentenced,convicted,
administrativa	administration,administrative,administative,
åtal	prosecution,
bin	bin,
dubbelt	double,
bil	car,
teknik	technique,technology,technic,
big	big,
kejsaren	emperor,the emperor,
avlidna	diseased,deceased,the perished,
af	of,of (old swedish),
möttes	met,
bit	piece,
indonesiska	indonesian,
planeterna	the planets,planets,the planet's,
rené	rene,rené,
grå	gray,grey,
kolonialtiden	the colonial times,colonial period,
angränsande	adjoining,adjacent,
möjlig	possible,
stränga	severe,
avsedda	aimed,for,intended,
tillstånd	state,to the dental,condition,
anatomi	anatomy,
google	google,
identisk	identical,
egyptiska	egyptian,
tolkningar	interpretations,interpretation,
back	reverse,
körberg	körberg,
historisk	historic,historical,
studerar	study,studies,
cocacola	coca cola,coca-cola,
lars	lars,
västergötland	västergötland,
flygplatser	airports,air ports,
måste	have to,must,
lasse	lasse,
integration	integration,
per	per,
pratar	talks,talking,talk,
självstyre	autonomy,self-governance,self-government,
saab	saab,
lösningen	the solution,solution,
därför	because,therefore,
nordamerika	north america,
resande	travelers,travelling,
vasaloppet	vasaloppet,
påven	the pope,paven,pope,
ockuperade	occupied,
britannica	britannica,
korta	short,
värmestrålningen	heat radiation,
uppfattningar	opinions,perceptions,
fallit	fallen,fall,
jimmy	jimmy,
grammy	grammy,
styrelse	government; direction,board,board of directors,
barcelonas	barcelona's,barcelona,
steven	steven,
ordnar	fix,decorations,arrange,
brita	brita,
paret	pair,the couple,parathyroid,
framträdde	appeared,emerged,
ökningen	increase,the increase,
dalar	valleys,
turkiska	turkey,turkish,
medvetande	consciousness,consciousnesses extensive,awareness,
lyssnar	listen,listens,
jaga	course,hunt,chase,
serie	comic; row; succession; serial,cartoon,series,
konsul	consulting,consul,
bostäder	residences,housing,
torsten	torsten,
oktober	october,
skillnaden	the difference,
ledningen	conduit,the lead,
mångfald	diversity,variety,
planet	planet,
smycken	jewlery,jewellery,
sultanen	sultan,
planer	plans,
amfetamin	amphetamine,
skillnader	differences,
reggaen	reggae,the reggae,
jordbävningen	the earthquake,earthquake,
reidar	reidar,
titel	title,
expedition	caretaker,expidition,expedition,
förbjudna	forbidden,prohibited,
hjärnans	the brain's,brain,
tropiskt	tropical,
tropiska	tropical,tropic,
materia	matter,materia,
tyskland	germany,
eller	or,
voltaire	voltaire,
familjer	families,
årstiderna	seasons,the seasons,
familjen	the family,family,
betalar	paying,pay,
makedonien	macedonia,
anser	believes,view,
anses	be,deemed; regarded,
maos	maos,mao's,mao,
lena	lena,
utvecklade	developed,oral,
länders	countrie's,countries',countries,
samla	collecting,collect,gather,
mutationer	mutations,
nådde	reached,
ritualer	rituals,
storkors	the grand cross,
talades	spoken,spoken (of),spoke,
regionala	regional,
sambandet	the connection,connection,relation,
dramatiker	playwright,dramatist,dramatists,
judisk	jewish,jew,
sorg	grief,sad,
regionalt	regional,regionally,
at	at,
flod	basin,river,
uppgår	is,shall amount,
jason	jason,
stänga	close,off,
stred	fought,
uran	uranium,
frankrike	france,
förut	requires,before,
sigmund	sigmund,
övergav	abandoned,
intensivt	intensive,hard,
privat	private,
lilla	small,
tillämpningar	applications,implementations,situations,
landslaget	the national team,team,
betrakta	view; regard,view,
sydafrikanska	south african,african,
sahlin	sahlin,
konsten	art,the art,
intensiva	intensive,intense,
kollaps	collapse,
atlas	atlas,
graven	the grave,grave,
passiv	passive,
luleå	luleå,
kampanjen	campaign,
plikt	duty,
turkiets	turkey's,turkeys,
annika	annika,
tjänade	earning,earned,
varnade	warned,
utgjordes	was,make up,comprised; consisted,
nonsporting	non sporting,
svts	svt,svts,
tävlingar	competitions,contests,
exemplet	the example,example,
knight	knight,
joel	joel,
samman	together,
slutade	quit,ending,
madeira	madeira,
warszawa	warzaw,warsaw,
endast	only,merely,
joey	joey,
tunnlar	tunnels,
störtades	overthrew,overthrown,was overthrown,
överhöghet	supremacy,suzeranity,sovereignty,
utbredda	widespread,spread,
vanligaste	frequent,most common,
cellen	cell,the cell,
påsken	easter,
earth	earth,
carlo	carlo,
depression	depression,
sträcker	stretches,extend,
går	is,goes,
chicago	chicago,
spåras	trace,
tillkomst	origin,established,advent,
senare	latterly; later,later,
sauron	sauron,
placering	position,placement,
rankning	ranking,rating,
analsex	anal sex,
och	and,
kyrka	church,
öar	islets,islands,
extremt	extremely,extreme,
ordförande	chairman,
luis	luis,
extrema	extreme,
isländska	icelandic,
befolkningstäthet	population density,the population density,
populäraste	rated,most popular,
störning	noise,
honom	his,him,
svårigheter	difficulties,hardships,
medeltid	medieval,the medieval times,
turkar	turks,
alaska	alaska,
lagts	added,
katolicismen	catholisism,catholicism,
lagförslag	bill,lagforslag,
miljard	billion,one billion,
honor	ära,female,
färgade	colored,
existens	existence,
protokoll	protocol,
uppnår	achieve,reaches,
uppnås	obtained,is achieved,
talare	speakers,speaker,spoke,
privata	private,
stundom	sometimes,somtimes,
når	reach,reaches,
nås	reached,is reached,
filippinerna	filipinos,the philippines,
betraktas	considered,
betraktar	regard,sees,
ovan	above,
lima	lima,
somrarna	the summers,summers,
skivbolag	record label,record company,
kinesisk	chinese,
skotsk	scottish,
chi	chi,
gruppspelet	group stage,groupplay,group play,
fånga	capture,capturing,
nobel	nobel,
döpt	named,baptized,
söder	south,
nytta	from,good,useful,
geografisk	geographic,geographical,spatial,
titanics	titanic's,titanic,
konkurrens	competition,
prinsen	prince,the prince,
platser	points,places,
förstå	understand,understandable,first,
utropade	exclaimed,cried out,
bakterier	bacteria,
självständighet	independance,independence,
avsikten	intention,purpose,
iii	iii,
platsen	the place,place,site,
ansvaret	responsibility,the responsiblity,
britney	britney,
f	f,
tunnel	tunnel,
gabriel	gabriel,
påbörjas	start,begin,starts,
halt	content,stop; level,stop,
baserad	based,
kedja	chain,
kategorisvenska	category: swedish,
baseras	based,bases,based on,
baserar	base,based,
baserat	based,
kyrkan	the church,church,
väldet	empire,violence,the rule,
indianerna	the indians,indians,
titlar	titles,
do	do,
mozarts	mozart's,mozart,
cecilia	cecilia,
fett	fat,
framtida	future,
internationellt	international,internationally,
lanserade	introduced,launched,
internationella	international,
tjänst	service,
vilhelm	vilhelm,
revs	described,was demolished,
böckerna	books,
rousseau	rousseau,
riktig	real,
klar	clear,done,
trycktes	was published,printed,
föddes	was born,born,
herrlandskamper	herrlandskamper,men's international contest,men's international contests,
brändes	burned,burnt,
spannmål	grain,cereals,
förbundskapten	manager,coach,
klan	clan,
gammal	old,
terrier	terriers,terrier,
siv	siv,
finländska	finish,finnish,
rådhus	town hall,courthouse,
dryck	beverage,drink,drinks,
förekommit	occured,occurred,
billboardlistan	billboard list,bilboardlist,
grannar	neighbors,neighbours,
registrerade	data,noted,
olyckan	incident,the accident,
alltjämt	remains,
bilbo	bilbo,
omslaget	cover,the cover,
dy	younger,
halvklotet	hemisphere,
strid	conflict,fight,
georg	georgian,georg,
innebär	mean,means,
industrier	industries,
le	smile,le,
människor	human,people,
la	la,
variationer	variations,
berget	mount,the mountain,
föreställer	picture,depicts,pictures,
tillägg	addition,appendix,
eus	eu,
dag	dag,day,
spektrum	spectra,spectrum,
utfärdade	issued,
slags	kind,type,
dam	dam,lady,
dan	dan,
valet	selection,the election,
avslöjar	reveals,
tillkommit	been,accured,
periodiska	periodic,
das	das,
sammanhanget	connection,context,
installera	installing,install,
day	day,
kontinuerligt	continuous,continous,
beslut	decision,
morris	morris,
newtons	newton,newton's,
syftade	alluded to,aiming,aimed,
spridningen	spread,proliferation,the spread,
lysande	brilliant,illuminating,
engelskspråkiga	english-speaking,the english language,
juridisk	legal,
krita	chalk,
humanism	humanistic,humanism,
pitts	pitts,
kristiansson	kristiansen,kristiansson,
dokumentär	documentary,
inspirerade	inspired,
segern	the victory,victory,
marley	marley,bob marley = singer,
arbetskraft	workforce,labor,
fattigdomen	poverty,
nödvändiga	necessary,essential,
matt	matt,dull,
jerusalem	jerusalem,
mats	mat's,attention,
kärnan	core,the core,
nödvändigt	neccessary,necessary,
deras	their,
red	eds,
återta	retake,regain,reclaim,
filmatiseringen	film version,
roterande	rotating,
frank	franks,
webbplats	website,site,
franz	franz,
odlas	cultured,
arbetare	workers,
ronald	ronald,
längre	longer,
josé	jose,
fart	off,speed,
efterträddes	succeeded,
medelhavsområdet	mediterranean,the mediterranean region,the mediterranean area,
referenser	references,
farbror	uncle,
striderna	the battles,fighting,
nivå	niva,level,
south	south,
liberaler	liberals,
klassisk	classical,classic,
genomgår	undergoes,undergoing,
pga	because of (short of "på grund av"),due,
uppges	reported,
uppger	states,state,
innehålla	include,contain,
insikt	insight,recognition,
levnadsstandarden	the standard of living,living standard,standard of living,
fruktade	feared,
omständigheter	event,circumstances,
veckan	weeks,the week,
leder	leads,leading (to),lead,
utlopp	outflow,outlet,
energikällor	energy resources,energy sources,sources of energy,
kantonerna	the cantons,cantons,
förklara	explain,declaring,
maidens	maidens,
leden	hinge,lines,the route,
palestina	palestine,
demonstrationer	demonstrations,
bundna	tied,bonded,bound,
noterade	note,noted,
stället	instead,the place,
ställer	running; causing,set,run (in election),
innehade	held,possessed,
firades	celebrated,was,was celebrated,
pågående	current,ongoing,
sjögren	sjögren,
ledamöter	commissioners,members,
släkten	genera,the family,
ställen	spots; places,places,
bevarats	protected,preserved,
beskrivningen	description,
domaren	judge,the judge,
matematisk	mathematical,mathematic,
inne	inside,in,
sweden	sweden,
kvalificerade	qualifying,
universum	universe,
mälaren	mälaren,
premiär	prime,premiere,
havs	at sea,sea,
aristoteles	aristoteles,aristotle,
tids	time,
operativsystem	operative systems,os,operating system,
följd	following,effect,
älgar	moose,
följa	following,follow,
basist	bassist,
uganda	uganda,
idag	today,
rådande	current,prevalent,
följt	followed,
följs	followed,
låt	let,song,
mil	mile,swedish miles,mil,
min	my,
mia	mia,
fötter	feet,on its feet,
kroppar	cells,bodies,
tidningar	press,magazines,
mig	me,
mix	mix,
låg	low,
experter	experts,
besättningen	crew,
lån	loan,
konstverk	work of art,artworks,artwork,
konkurrerande	competing,
kommunikationer	communications,
resurser	resources,
resultatet	the result,result,
dinosaurier	dinosaurs,
varandras	each other's,each others,each other,
missionärer	missioners,missioner,missionaries,
resultaten	the results,results,
sedan	then,since,
sist	finally,last,
efternamn	last name,lastname,surname,
liknade	looked like,similar,
stranden	shore,the beach,
upprustning	renovation,
irakkriget	iraq war,
republikanska	republican,
rörelsens	movements,operating,movement,
milano	milano,
deuterium	deuterium,
tidskrift	newspaper,magazine,
capita	capita,
styrke	strength,been,
definiera	defining,define,
viktigaste	most important,
styrka	strength,power,
utgångspunkt	starting point,point of departure,
obelix	obelix,
text	text,
komplicerad	complex,complicated,
existerande	current,existing,
hamlet	hamlet,
inhemsk	domestic,native,
ugglas	owl,ugglas,
fungerade	thought,working,
kurfursten	elector,
rumänska	romanian,
järnvägen	railroad,rail,
euroområdet	eurozone,euro area,convergence report,
rytmiska	rhythmic,more rhythmic,
satan	satan,
shahen	the shah,shah,
säker	items,safe,safety,
bryssel	brussels,
organiska	organic,
snitt	on average,average,
arean	the area,the space,area,
förändrades	changed,
buddhismen	buddhism,buddism,buddhismen,
överlägset	far,superior,
förstår	understand,forstar,
regimen	regime,
studenterna	students,the students,
uppehåll	residence,pause,hiatus,
richards	richards,
från	from,
vinsten	the win,gain,
organ	body,agency,organ,
županija	country,
nazitysklands	nazi germany's,nazi germany,
vinster	profit,gains,
majoriteten	the majority,
lyckade	successful,
byggdes	was,was built,
ronaldo	ronaldo,
militärer	military,soldiers,
krävdes	were required,
national	national,
svenska	swedish,
eleonora	eleonora,
kapitalet	the capital,capital,
svenskt	swedish,
först	first,
bön	nests,prayer,
debutalbumet	the debut-album,debut album,
reform	reform,
redan	already,has already,
konverterade	converted,
seder	subsequently,custom,
bruno	bruno,
carlsson	carlsson,
avslutades	closed,ended; concluded,concludes,
vänta	(have to) wait; expect,wait,
bör	live,should,
terräng	terrain,off,
ordentligt	proper,properly,firmly,
översikt	overview,over term,
koncept	concept,
industrialisering	industrialization,
tobias	tobias,
uppskattade	estimated,appreciated,
listan	the list,
hårdare	harder,more severely,tougher,
säkerheten	the security,safety,
översättas	translated,be translated,translated (to),
viktigare	important,more important,
läsning	read,reading,
hämtade	taken,brought,
buddhas	buddha's,buddhas,
empathy	empathy,
miniatyr|karta	thumbnail map,miniature|map,
återförening	reunion,
litteratur	literature,litterature,
aktuellt	current,relevant,
kommunicerar	communicates,
kröntes	been crowned,crowned,
aktuella	current,
kommendör	commandor,commander,
förekomst	presence,
sachsen	sachsen,saxony,
fester	celebrations,parties,
inneburit	meant,resulted,
befogenhet	warrant,authorization,authority,
utsågs	was,appointed,was appointed,
medicinsk	medical,
elektroner	electron,electrons,
news	news,
ad	ad,
västmakterna	western powers,
tunisien	tunisia,
grupperingar	groupings,groups,grouping,
slippa	avoid,
gaza	gaza,
igen	again,back,recognize,
define	define,
asteroider	astroids,asteroids,
genomsnittlig	average,
stationen	station,
stationer	stations,
lärjungar	disciple,disciples,
deep	deep,
uppmärksammat	attention,noticed,
an	an,
napoleon	napoleon,
augusti	august,
bruket	use,the use,
kraftiga	strong,powerful,
stalin	stalin,
ar	is,
ocheller	and/or,
betraktade	considered,watched,
externa	external,
palats	palaces,palace,
tagits	taken,
flyktingar	refugees,
betalade	payed,paid,
fördrag	agreement,treaty,
vistelse	visit,stay,
prosa	prose,
videon	the video,video,
händelserna	the events,events,the happenings,
administration	administration,
lämnade	did,left,
wolfgang	wolfgang,
blodtrycket	the blood pressure,blood pressure,
sångerna	song are,the songs,
omedelbart	immediately,immediate,
heinrich	heinrich,
hinduismen	hinduism,up,
kallad	known as the,know as,called,
kontrollera	control,controlling,
framförallt	above all,in particular; above all,
kallat	called,
kallas	called,
kallar	call,calls,
center	center,
öde	fate,
seth	seth,
antonio	antonio,
sett	seen,except,
hoppas	hope,
omgångar	in turns; periods; mandates,cycles,
svensk	swedish,
undvika	prevent,avoid,
position	position,
deltar	part,participates,
innehåll	content,contents,
stores	great,the great's,the great,
kontaktade	contacted,
passade	suiting,suited,fit; suited,
mystiska	mysterious,mystical,
wagner	wagner,
misshandel	assault,abuse,
grekiskans	the greek's,greek,
flertal	several,majority group,
vanligt	usual,normal,
hamburg	hamburger,hamburg,
kampf	on,kampf,
liverpools	liverpool's,liverpools,
reformer	reformers,reforms,
anhöriga	relatives,kin,
lake	lake,
mentala	mental,mentala,
landområden	land,land areas,
streck	bar,
match	game,match,
förnuft	common sense,reason,
uppmärksamhet	attention,attantion,
uppträder	appears,performs,occur,
dubai	dubai,
demens	dementia,
innehöll	containing,include,
chrusjtjov	khrushchev,chrusjtjov,
viruset	virus,
likt	like,
journalist	journalist,
works	works,
uppträda	occur,appear,act,
gudomlig	divine,
albumets	album,album's,
starkaste	strongest,the strongest,
insats	contribution,intermediate,stake,
etablerades	established,was established,
minsta	minimum,
est	est,
joachim	joachim,
katarina	katarina,
löser	solve,solves,
skildrar	depicts,describes,portrays,
kategorifiktiva	category fictitious,
gisslan	hostage,hostages,
internationalen	international,
definitionen	definition,the definition,
nattetid	overnight,
definitioner	definitions,
starkare	strong,stronger,
leopold	leopold,
arterna	the species,species,
nordkorea	north korea,north koreans,
socker	sugar,
ärkebiskopen	archbishop,
glada	happy,
mäktigaste	powerful,most powerful,
slutgiltiga	final,
andel	percentage,share,
anden	the holy spirit,spirit,
folkräkningen	census,
värd	host,worth,
alexanders	alexanders,alexander's,
förstärka	strengthen,enhance,
kapital	capital,
omgiven	surrounded,
potatis	potato,
monarken	the monarch,monarch,
chris	chris,
australiska	australian,
ljusare	brighter,lighter,
föredrar	prefer,preferred,
vimmerby	vimmerby,
hatar	hate,hates,
ridge	ridge,
densamma	the same,same,
skog	wood,forest,
kuben	cube,the cube,
möjliggjorde	made possible,enabled,allowed,
föga	little,hardly; little,
flyg	flight,airforce,air,
kärnor	core,cores,
kväll	evening,
klockan	clock,o'clock,
civilbefolkningen	civilian population,the civilian population,civilians,
ryssarna	the russians,russians,
brand	fire,
bröder	brothers,
ersättning	pay,replacement,
flygvapnet	air force,the airforce,
kraft	force,power,
bud	bid,bids,message,
nöjd	content,
vetenskap	science,
utrymme	space,
arbetsgivaren	employer,
individens	individual's,the individual's,
australiens	australia,australia's,
nedre	lower,bottom,
kaffe	coffee,
minuter	minutes,
vänstra	left-hand,left,
hästens	horses,horse's,horse,
circus	circus,
paraguay	paraguay,
tolkningen	interpretetation,interpretation,
omloppsbanor	orbits,orbit,
autism	autism,
betydande	important,significant,
kommuner	municipalities,local,counties,
manlig	male,manly,
identitet	identity,
särskilda	specific,special,
proteinet	protein,the protein,
proteiner	proteins,
einsteins	einstein,once a,einsteins,
uppfattar	sees,percieves,interpret,
picchu	picchu,
stimulans	stimulation,stimulating,
betonade	emphasized,
uppfattas	be perceived,perceived,are regarded,
försämrades	worsened,worsening,decreased,
uppfatta	apprehend,perceived,perceive,
sjön	lake,
tämligen	rather,fairly,tamil again,
astronomi	astronomy,
variation	diversity,variety,
koncentrationsläger	concentration,concentration camp,concentration camps; kz-camps,
akademisk	academical,academic,
ärkebiskop	archbishop,
cirkel	circular,
philips	philips,
fakta	facts,fact,
winnerbäck	winnerbäck,winnerback,
baker	baker,
svag	weak,
uppfattningen	comprehension,view,
framför	in front of,particularly,above,
förbundet	the union,association,
okänd	unknown,
nelson	nelson,
mäktiga	powerful,
brottslingar	criminals,
nederländerna	the netherlands,netherlands,
båt	boat,
resor	travels,travel,
påsk	easter,
arkitekt	architect,
antisemitiska	antisemetic,anti-semitic,antisemitic,
ozzy	ozzy,
granskning	review,
anfallet	the attack,attack,
upphör	end,
paris	paris,
tillväxten	growth,
deltagit	part,participated,
kapacitet	the capacity,capacity,
under	during,for,under,
läge	mode,location,
svårare	harder,difficult,
nordost	north east,northeast,the northeast,
pommern	pommern,pomerania,
ägande	owning,ownership,
socialdemokrater	social democrats,
jack	jack,
invånare	resident (-s),inhabitants,
evert	everted,evert,
kammare	chamber,
tagit	taken,received,
school	school,
utmärks	are characterized,characterized,
utmärkt	excellently,excellent; superb; marked by; characterized by,excellent,
öppna	open,
plural	plural,
venus	venus,
matematik	mathematic,mathematics,
verklig	real,
reklam	advertising,advertisement,
parten	party,
markerar	selects,marks,
kropp	body,
bönderna	the farmers,farmers,
manus	script,
läget	position,location,
indierna	the indians,indians,
läger	camps,camp,
stridigheter	oppositions,strife,
aktivt	active,actively,
drivande	drive,driving,
ebba	die,ebba,
notera	note,
liberty	liberty,
aktiva	active,
zink	zinc,
kub	cube,
disney	disney,
egyptens	egypt,egypts,egypt's,
språken	languages,park,
zach	zach,
prata	talk,
flera	many,multiple,
medelhavsklimat	mediterranean climate,
utredning	study,investigation,
beck	beck,pitch,
parlamentariska	parliamentary,the parliamentary,
preparat	substance,preparations,compound,
studio	studio,
rysk	russian,
sommartid	summer-time,summer,during summer,
komplex	complex,komplex,
studie	study,
språket	language,
forum	forum,
lagras	stored,
ty	for,
precis	precisely,exactly; precisely,just,
proportioner	proportions,
svante	svante,
gällande	current,regarding,
koloniserades	is colonized,colonized,
upptäckter	discoveries,discovery,
upptäcktes	discovered,(was) discovered,
julie	julie,
erektion	erection,
julia	julia,
övers	transl,translation,
nazistiska	nazi,
misslyckats	failed,
upptäckten	the discovery,discovery,
försvarsmakt	armed forces,
eftervärlden	posterity,the world,
volym	volume,
mattias	mattias,
klassas	classified,
vinst	profit,win,
miniatyr|px|en	miniature,
konserterna	the concerts,concerts,
västtyskland	västttyskland,west germany,
skicka	send,
behandlingar	treatments,
belägg	coating,evidence,
återstående	remaining,
muse	muse,
övertala	convince,persuade,
ludvig	louis,ludvig,
ansökte	applied,
världsarv	world heritage,
fermentering	fermentation,
rörelse	movement,
belgiens	belgium,belgium's,
igelkottens	the hedgehog's,hedgehog,
henri	henri - it's a name,henri,
mm	millimeter,etc.,
arméns	the army's,arm,army's,
lukas	luke,lukas,
antiken	the ancient world,antiquity,
ms	motor ship,
mr	herr,mr,
johanssons	johanssons,johansson,
ernest	ernest,
avstå	desist,non,refrain,
utgick	started,was deleted,
partiets	the party's,parties,
ghana	ghana,
sträckan	distance,the distance,
utlöste	triggered,
persien	persia,
trädgård	garden,
florida	florida,
genomfördes	completed,was,was carried out,
fröken	miss,
ena	one,
end	end,
smält	melted,
iiis	iii's,3's,
väpnade	armed,
ens	even,one's,
gata	street,
elektriskt	electric,
elizabeth	elizabeth,
beskrev	depicted,described,
målen	cases,goals,
förståelse	understanding,
mest	most,mostly,
västvärlden	west,western world,
målet	target,the target,
miniatyr|px|ett	miniature,
elektriska	electrical,
frågade	asked,
 cm	centimeters,cm,
nagasaki	nagasaki,
kategorier	categories,
kubanska	cuban,
galilei	galilei,
beteenden	behavior,
kontrollen	control,the control,
existera	exist,
beskrivit	described,
praxis	practice,
arbetar	work,works,
kejsare	emperor,
kampen	the struggle,the fight,fight,
over	over,
arresterades	was arrested,
vitt	white,widely,
london	london,
synonymt	synonymous,synonymously,
frivillig	optional,
vita	white,
expansion	expansion,
bibelns	the bibel's,the bible's,bible,
brinner	on fire,burns,burn,
evans	evans,
imf	imf,
edith	edith,
nytt	new,
statschef	head of state,
dött	dead,died,
blott	merely,only,mere,
historiens	historys,history's,
dem	those,
senast	last (time),last,
produktion	production,
upptagen	included,busy,occupied,
avskaffandet	elimination,abolition,abolishment,
ansvarar	charge,responsible,
alex	alex,
jämförelser	comparison,
detroit	detroit,
bunny	bunny,
ställdes	was positioned,prepared,
newport	newport,
storlek	size,
ursprungligen	initially,originally,
växter	plants,
önskemål	desire,requests,demands,
gymnasium	high school,
group	group,
bra	good,
dessförinnan	before (that),before,
träffade	met,
innehållande	containing,including,
platina	platinum,
näst	second,second (to),
nio	nine,
medelålder	middle age,mean age,
behövs	required,is needed,
god	good,
receptorer	receptors,
användningen	use,the use,
ammoniak	ammonia,
hemland	homeland,
riktning	direction,
danmarks	denmarks,denmark's,
paulus	paulus,paul,
got	got,
behöva	need,
independence	independence,
smala	narrow,
bröderna	brothers,the brothers,
icke	non,none,
herman	herman,
värnplikt	military service,
kandidat	candidate,
fred	peace,
statsöverhuvud	head of state,
undervisade	taught,
samlade	collected,
inom	within,in,
drygt	good,approximately,
statsministern	the prime minister,prime minister,head of state,
studera	study,
tolerans	tolerance,
bredvid	beside,next to,
vetenskapliga	scientific,
hjälpte	helped,
befolkade	inhabitated,populated,
vetenskapligt	scientifically,scientific,
transporterar	carrying,transports,
transporteras	is transported,transported,
nyheter	news,
säsong	season,
museet	the museum,museum,
museer	museums,musser,
föreslagits	suggested,was suggested,
nhl	nhl,
institutioner	institutions,
rikaste	the richest,richest,
tillåts	is allowed,allowed,
yngsta	youngest,
sexuella	sexual,
nyheten	news,
mercury	mercury,
vikingar	vikings,
tor	thu,thor,
yngste	youngest,
punkten	the point,point,
à	à,river,
konventionen	the convention,convention,
merkurius	mercury,
å	on,river,of the,
konventioner	conventions,
ton	tonne,tone,
punkter	points,seq,
tom	tom,
uppkommit	generated,arisen,
tog	was,took,
fördes	sea were entered,out,
adjektiv	adjective,adjectives,
ifrågasatts	is questioned,questioned,
livealbum	live album,
skildes	separated,was seperated,
meddelande	message,
rädsla	fear,
fördel	advantageously,advantage,
kulturarv	culture heritage,cultureheritage,cultural heritage,
territoriella	territorial,
dramer	dramas,plays,
slutsats	conclusion,
mjölk	milk,
uppmuntrade	encouragement,encouraged,
bridge	bridge,
rad	range,line,
nedgång	decline,decreases,fall,
flyttades	moved,
tänka	thinking,think,
rak	straight,linear,
somliga	some people,some,
störningar	interruptions,disorder,disorders,
växer	growing,grows,
ras	race,ras,
adhd	adhd,
övervikt	obesity,overweight,
tycks	appears,
tänkt	expected,supposed; intended,intended,
ray	ray,
industriellt	industrially,industrial,
hittats	found,
kvällen	the evening,evening,
situationer	situations,
jorden	the earth,earth,earth; earth; underground,
lanseringen	the release,launch,
användning	use,use; usage,
fartyg	vessel,ship; vessel,ship,
industriella	industrial,
academy	academy,
situationen	situation,the situation,
mekaniska	mechanical,
grundskolan	elementary school,
tvingas	forced,system,
skepp	vessel,ship,
elektricitet	electricity,
fralagen	fra law,fralegen,the fra law,
spelat	played,
framgångsrik	successful,
spelas	played,
tanzania	tanzania,
metal	metal,
sekt	sect,
metan	methane,
sjöar	lakes,parks,
inflytande	influence,power,
agnes	agnes,
utkanten	the outskirts,outskirts,
dyrare	more expensive,expensive,
idrott	sport,sports,
saga	saga,story,
järnvägarna	the railways,railways,
queen	drottning,
gränserna	borders,the borders,limits,
radio	radio,
höjdpunkt	highlight,climax,high point,
sagt	said,i have said,
radie	radius,
absolut	absolute,absolute; total,
skada	damage,
claude	claude,
florens	florence,florens,
vinna	win,
resterande	remainder,remaining,
ägare	owner,owners,
gods	domain,goods,
holländska	dutch,
abu	abu,
återstår	remains,remain,
andras	others,
länder	states,countries,
torah	torah,
kommunisterna	communists,communist,the communists,
guatemala	guatemala,
gogh	gogh,
haiti	haiti,
sträckor	distances,
ålder	age,
stadskärnan	town/city,city bear man,center,
taubes	taubes,
ändras	be changed,change,
ändrar	changing,changes,change,
ursäkt	excuse,apology,
ändrat	changed,modified,
lovat	promised,
publicerades	published,
tidningen	the newspaper,journal,paper,
utvisning	penalty,expulsion,
kroppen	body,the body,
sakta	slowly,
ockuperat	occupied,
fördomar	bias,prejudice,prejudices,
kristendomen	chritianity,christianity,
utformade	formed,designed,
behålla	container,keep,
mur	wall,
indoeuropeiska	indo-european,european,
brinnande	burning,
antikens	the ancient's,ancient,
populär	popular,
slottet	castle,the castle,
finger	finger,finder,
förstås	course,mean:,
allra	very,most,-most; most,
mun	mouth,oral,
herding	herding,
förhållande	in relation,ratio,(in) comparison (to),
ordnade	arranged,parent,
betonar	stress,emphasize,
maniska	manic,maniac,
seden	the seed,custom,
dödsorsaken	cause of death,
bildriksdagsval	image election,
nummer	number,
store	great,
börje	börje,borje,
kreativitet	creativity,
autonomi	autonomy,
anfall	attack,
verka	seem,operate,appear,
lösningsmedel	solvent,
läggs	is,put before; submitted; put,lay,
farliga	dangerous,
allierades	allied's,allied,
begränsade	restricted,limiting,
förbränning	combustion,incineration,
avgöra	determine,decide,
lägga	put,add,lay,
grupper	groups,
hitler	hitler,
solljus	sun light,sunlight,
skapades	generated,created,
rumänien	romania,
grundaren	the founder,founder,
strävhårig	hispid,wirehaired,
aktiv	active,
hastighet	speed,
diktatorn	the dictator,dictator,
homosexuell	homosexual,
skalan	scale,
öster	east,
modernare	mor modern,more modern,
anspråk	claims,claim,
spritt	spread,
börja	start,
drömmar	dreams,
invasionen	invasion,the invasion,
älgen	elk; moose,moose,
n	n,
petrus	petrus,
schizofreni	schizophrenia,
depp	depp,
förståelsen	the understanding,
claes	claes,
della	della,
nationer	nations,
född	born,
darwins	darwin,darwins,
därigenom	by which,thus,thereby,
vojvodskap	voivodships,voivodeship,
brott	breach,crimes,crime,
anlände	arrived,
känsliga	susceptible,1st&2nd: fragile 3rd: sensitive,bilge accordance,
nationen	the nation,
kartan	the map,map,
vanföreställningar	delusions,
varefter	whereafter,
ekonomin	the economy,economy,
väljs	selected,elect,
ernman	ernman,
äger	owns,
rna	rna,
pekar	points,pointer,pointing,
erhållit	obtained,acquired,received,
ökade	increased,
ersatte	substituting,replaced,
pekat	pointed,identified,
negativ	negative,
welsh	welsh,
hundra	hundred,one hundred,
formatet	the format,size,format,
ersatts	replaced,(has been) replaced,
återvände	returned,returning,
återvända	return,
uppsving	boost,
gudom	deity,
dylan	dylan,
charlie	charlie,
spelad	played,
tillkännagav	announced,
svavel	sulfur,sulphur,
kemikalier	chemicals,
fattigare	poorer,
louisiana	louisiana,
jean	jean,
motsatt	opposite,
motsats	contrary,
spelar	gaming,
mytologin	mythology,
kraftigt	heavily,
järn	iron,kon,
ämnen	agents,substances,
mängd	volume,amount,laden,
graden	rate,the degree,degree,
europaparlamentet	european-parliament,the european parliament,european parliament,
grader	degrees,
engelskans	english,
utföras	be,performed,
kolväten	hydrocarbons,the hydrocarbon,
kalifornien	california,
använt	using,used,
värnpliktiga	conscripted,inductees,
gavs	was,gave,
belagt	coated,
eld	fire,
reglera	expell,controlling,
därefter	then,thereafter,
rätta	correct,come to grips; court; correct,
regionerna	regions,
enlighet	union,according (to),according,
 au	au,
benämning	term,name,title,
donau	the danube,danube,donau,
ämnet	substance,subject,
tillgänglig	available,provided,
protesterade	protested,
auktoritet	authority,
omvärlden	world,surrounding world,outside world,
gift	married,
såväl	both,as well as,
ladda	load,
modersmål	native language,mother tongue,
bosnienhercegovina	bosnia-hercegovina,
specifik	specific,
tillåtna	allowed,
fotbollen	soccer,football,
hund	dog,
gifter	marries,toxins,
lagstiftningen	law-making,legislation,
varianterna	variants,the diversities,
hanhon	he/she,male-female,
hushåll	household,
besöka	visit,
jennifer	jennifer,
malaysia	malaysia,
donald	donald,
besökt	visited,
saturnus	saturn,saturnus,
skapa	create,creating,
estetik	esthetics,aesthetics,
ultraviolett	ultraviolet,
totalt	total,complete,wholly,
användare	users,
gösta	gösta,gosta,
icd	icd,
diktatur	dictator,dictatorship,
utse	appoint,name,
tjorven	tjorven,
totala	total,
karaktäriseras	characterizes,is characterised,is charactarized,
elitserien	elite series,elitserien,
monoteism	monotheism,
ishockeyspelare	hockey player,ice hockey player,hockey players,
tillbringar	spends,spend,
män	males,men,
spelare	player,
hotellet	the hotel,hotel,
meyer	meyer,
census	census,
titeln	the title,title,
tvingades	forced,had,
systrar	sisters,
omgången	round,
plus	plus,
analytisk	analytical,
internationell	international,
hår	hair,
tydliga	clear,obvious,
kvarstår	remains,
primitiva	primitive,
civil	civil,civilian,
menade	meant,said,
systemet	the system,system,
tydligt	clear,obvious,
isberg	ice berg,iceberg,
sinne	mind,
anorexia	anorexia,
oförmåga	inability,failure,incapacity,
omges	surrounded,
omger	surrounds,surrounding,surrounding the,
lagt	laid,added,
kjell	kjell,
sicilien	sicily,
anderson	anderson,
kronprinsessan	crown princess,
metabolism	metabolism,
wittenberg	wittenberg,
dialekterna	dialects,
fadern	the father,
skulden	the debt,the guilt,
barrett	barett,barrett,
fängelsestraff	imprisonment,prison,
italien	italy,
skulder	debts,liabilities,debt,
finns	is,exist,there is,
eventuell	any,
fusionen	merger,the fusion,
säkerhet	safety; security,security,
amerikanerna	americans,the americans,
värvade	recruited,referred,
tillika	also,well,
araber	arabs,
behandla	treatment,
trio	trio,
bildt	bildt,
everest	everest,
bilda	form,
läsa	read,
tronen	throne,the throne,
generna	genes,the genes,
förbud	ban,prohibiting,prohibition,
liberalism	liberalism,
tätorten	conurbation,agglomeration,
ni	you,
margareta	margareta,
no	no.,
tillverkade	manufactured,made,
when	when,
nf	nf,
finna	found,
ny	new,
tio	ten,
lösas	solved,
nr	no.,number,no,
tätorter	urban,conurbation,cities,
nu	now,
picture	picture,
phoenix	phoenix,
sätts	is,turned (on),is placed,
miscellaneous	miscellaneous,
gäster	guests,
tunna	thin,
massakern	massacre,
sätta	insert,set,
kronprins	crown prince,
väckte	awakened,aroused,
beroendeframkallande	addictive,
vietnam	vietnam,
cellens	the cell's,cell's,the cells,
rom	rome,rom,
ron	ron,
rob	rob,
rod	rod,
dvärg	dwarf,
roy	roy,
koreanska	korean,
udda	odd,
minska	reducing,reduce,
laura	laura,
mottagarens	the reciever,the receivers,the receiver's,
konstitutionell	constitutional,
bär	carryng,berries,here,
tanke	light,in light of,
federation	federation,
även	even,also,
läns	county,county's,
varvid	in which,
underhållning	entertainment,
flytt	escaped,move,fled,
forna	former,previous,
metod	method,
inlärning	learning,
brother	brother,
christmas	christmas,
olyckor	accidents,
lever	living,live,liver,
länkar	links,
församling	congregation,assembly,
införandet	introduction,the introduction,
trend	trend,
stilar	styles,
kategorirock	category:rock,category rock,
linda	winding,linda,
colin	colin,
svartån	svartån (black stream),svartån,
förorter	suburbs,
port	gate,port,
uppgifterna	the information,data,
ifråga	with regards to,in question,challenged,
poesi	poetry,
agnosticism	agnosticism,
miniatyr	miniature,thumbnail,
ögat	eye,
cykel	bicycle,cycle,
månaderna	months,
angelina	angelina,
gräs	grass,
gravitation	gravitation,gravity,
kamp	struggle,fight,
vindkraftverk	wind power station,wind turbine,
enkla	simple,single,
metaller	metals,
eiffeltornet	the eiffel tower,
jord	soil,earth,
turister	tourists,
dublin	dublin,
sina	their,his,
införts	been inserted,introduced,
lokal	local,
ankomst	arrival,
filmen	the movie,film,
tilltagande	increasing,
rafael	rafael,rafel,
bevara	preserve,preserving,
luften	air,
sikt	term,run,
etablera	establish,up,
trummor	drums,
bolaget	company,the company,
ungerska	hungarian,
russell	russell,rusell,
undan	away (from),escape,
utropades	proclaimed,was proclaimed,
samfundet	the communion,association,
lp	lp,
anda	spirit,
inblandade	involved,
andy	andy,
kurder	kurds,
australian	australian,
turné	tour,
crüe	crüe,
uppskattningar	estimates,
typerna	the types,types,
staten	state,
kär	in love,
övergå	transition,transend,
palestinsk	palestinian,
årets	the year's,year,
efterhand	post,hindsight,
piano	piano,
styras	guided,controlled,steered,
drabbades	affected,where hit by,afflicted,
läkemedel	drugs,medicine,
musikaliska	musical,
rådgivare	counsellor,advisor,
valla	wax,valla,herd,
jude	dude,jew,
allvarlig	serious,
judy	judy,
humle	hops,hop,
generell	general,
karibiska	caribbean,
musikaliskt	musically talented,musical,musically,
anpassat	adapted,
uppväxt	growing up,
bönorna	bean,beans,
bära	carry,mean,
dokumenterade	documented,
utdelades	distributed,awarded,
hemligt	secret,
annorlunda	different,otherwise,
hemliga	secret,
främja	further,promote,promoting,
swedish	swedish,
frivilligt	voluntarily,voluntary,
speglar	mirror,mirrors,
avrättning	execution,
frivilliga	volunteers,optional,voluntary,
andlig	spiritual,spirtual,
stöter	thrust,run,
simning	swimming,
regeln	the rule,rule,
muslimerna	muslims,the muslims,
inriktad	focused on,oriented,intent,
etablerat	established,
tvserien	tv series,the tv show,television program,
levt	survived,
fascism	fascism,
sydliga	southern,
familjens	the familys,family,
flög	fly,flew,
fenomen	phenomena,phenomenon,phenomenazaqq,
leva	live,
utrikespolitiska	foreign policy,foreign political,
väntan	awaiting,waiting,wait,
marknad	market,
kroniska	chronic,
beror	is,
stridande	conflict,fighting,warring,
japanska	japanese,
väntat	expected,
väntas	expected,
väntar	waiting,expect,
faser	phase,phases,
orter	varieties,locations,
kartor	maps,
bushs	bush,bush's,
orten	resort,the suburb,
födelse	date,birth,
komplicerat	complex,complicated,
iberiska	iberian,
fasen	phase,
rapport	report,
böcker	useful downloads archive,books,
kämpade	fought,
välja	select,
wallace	wallace,
undervisningen	teaching,the education,
sätt	manner,way,
förespråkare	spokesman,proponent,
behandlingen	the treatment,the treament,treatment,
spelarna	players,
försvaret	repository,the defense,
tjänstemän	officers of,officals,officials,
marleys	marley's,marley,
passar	suitable,suits,
hergé	herge,hergé,
femte	fifth,
hamilton	hamilton,
karlsson	karlsson,
tredjedel	a third,third,
hotar	threatens,
term	term,
opera	opera,operator,
snabb	instant,
namn	name,
futharkens	futharkens,futhark,the futhark's,
viggo	viggo,
alternativ	alternative,
hotad	threatened,
färger	color,colors,
bildning	education,form,learning,
semifinal	semifinals,semi finals,
förhandlingarna	the negotiations,negotiations,
stående	standing,above,
valuta	currency,exchange,
hoppade	jumped,
die	die,
amerikansk	american,u.s.,
åsikt	opinion,
behandlar	treats,treat,
behandlas	treated,
upprepade	repeated,
accepterad	acceptable,
stortorget	stortorget,the main square,
årliga	annual,
profil	profile,
accepterar	accepts,accept,
accepterat	accepted,
kent	kent,
malta	malta,
brett	broad,
juldagen	christmas day,
zuckerberg	zuckerberg,
etanol	ethanol,
nått	reached,
hjalmar	hjalmar,
pjäs	piece,
soundtrack	soundtrack,
arbetet	work,the work,
händelse	event,handel,
traditionen	the tradition,tradition,
motion	motion,exercise,
traditioner	traditions,the traditions,
place	place,
någonsin	ever,
politiken	policy,the politics,
hemsida	website,homepage,
blood	blood,
origin	origin,
begår	commits,commit,
såldes	sold,
självbiografi	autobiography,selfbiografi,
centralamerika	central america,
george	george,
respekt	respected,respect,
given	given,
ian	ian,
vågor	waves,
skjuten	shot,
cullen	cullen,
bahamas	bahamas,
skjuter	shoots,slide,extend,
givet	granted,given,
hud	skin,
personlighetsstörningar	personality disorders,
spelats	recorded,been played,played,
webbplatser	webbsites,websites,
gia	gia,
användandet	usage,use,
grund	in the context: "på grund" = because of,because,
montenegro	montenergo,montenegro,
alan	alan,
kallade	called,
nobelkommittén	the nobel commitee,
hur	how,the,cage,
hus	house,housing,a house,
webbplatsen	webpage,the website,site,
population	population,
smeknamn	nickname,
modellen	model,the model,
balans	balance,
marinen	navy,marines,
löfte	promise,
genomsnittet	average,the average,
framställning	preparation,production,
landsting	county,county council,
modeller	models,
bildades	founded,formed,was formed,
hjärtat	heart,the heart,
rena	pure,
mottagare	recipient,receiver,
ana	feel,ana,
tiotusentals	tens of thousands,
kromosomerna	chromosomes,the chromosomes,
maten	the food,
mando	command,
rent	true,clean,
jordskorpan	earth's crust,earth crust,the earth's crust,
världen	world,the world,
avstånd	distance,
förste	chief,the first,first,
första	first,
ideal	ideals,ideal,
förhållandena	conditions,the conditions,
gustavs	gustavs,gustav,
kust	coastal,coast,
periodvis	periodically,
stjärnornas	stellar,the star's,
knutna	associated,attached,tied,
diskussioner	discussions,discussion,
falla	fall,
 miljoner	one million,millions,millon,
invånarna	inhabitants,inhabitatants; citizens',residents,
staterna	states,usa,
täckt	covered,coated,
täcks	covered,covers,
lisbet	lisbet,
elektromagnetisk	electromagnetic,
erkänner	admits,recognize,
stövare	beagle,hound,
täcka	cover,thank,
tron	faith,
ronaldinho	ronaldinho,
mänskligheten	humanity,
bernadotte	bernadotte,
isolering	isolation,
sjunka	decrease,descend,
tror	believe,think,
bandets	the bands,band,
gula	yellow,
tvprogram	tv program,tv-show,
guld	gold,
tidningarna	papers,
flydde	fled,
motivet	the motive,subject,
ovanligt	unusual,rare,
gult	yellow,
iväg	away,off,
ovanliga	unusual,rare,
analys	analysis,
berättelser	tales,stories,
webbkällor	websources,webbkällor,web sources,
larsson	larsson,
aktiviteten	the level of activity,activity,
grundandet	founding (of),founding,
tränaren	coach,the coach,
jazz	jazz,
administrativ	administrative,administration,
nedåt	down,downward,down; downwards,
väder	weather,
theta	theta,
forsberg	forsberg,
mörkt	dark,
tränade	trained,
dramat	drama,the drama,
umeå	umeå,
joker	joker,
republika	republic,
osäkert	insecure,unclear,uncertain,
baltikum	the baltics,baltics,
satte	put,put together,sat,
minnen	memories,memory,
beethoven	beethoven,
tekniska	technical,
inspelningen	recording,
uppdraget	task; assignment,assignment,
tekniskt	technical,
college	college,
stanley	stanley,
minnet	the memory,memory,
älg	elk,moose,
freden	the peace,peace,
federal	federal,
utbud	range,availibility,supply,
skett	done,happened,
önskade	desired,wished,
översättning	translation,
återigen	once again,yet again,aterigen,
intresserad	interested,
hämtat	collected,downloaded,taken,
konstnären	artists,the artist,artist,
mellan	between,
antagligen	ligands presumably,probably,presumably,
konstnärer	artists,
bekämpa	prevent,combat; fight,fight,
ruiner	ruins,
dödade	killed,
myter	myths,
högre	higher,
come	come,
summa	sum,total,
sydeuropa	south europe,southern europe,
region	region,
ordagrant	literally,literal,verbatim,
spindlar	spiders,
lenins	lenin,lenin's,
introducerades	introduced,
gjorde	did,
gjorda	made,done,
pakistan	pakistan,
utgåvor	editions,issues,
regler	rules,
period	period,
pop	pop,
fransk	french,france,
werner	werner,
statens	state,the government's,
utformning	layout,shape,formation,
hävda	claim,asserting,
poe	poe,
skånska	scanian dialect,scanian,skånska,
howard	howard,
folken	the peoples,people,peoples,
strikta	strict,
förekomsten	existence,presence,
dagarna	the days,day,
musikstil	music still,music,music style,
folket	the people,people,
invaderade	invaded,
anderna	andes,the andes,
sändebud	messenger,envoy,
andres	andres,other's,
stadshus	city hall; town hall,town hall,
tjänster	services,
kapitulation	surrender,capitulation,
tiger	tiger,silent,
övrig	other,
minister	minister,
andré	andre,
kaos	chaos,
andrea	andrea,
champions	champions,
hughes	hughes,
användes	was used,used,
riktade	targeted,
mount	mount,
influenser	influence,influences,
cash	cash,
arnold	arnold,
spreds	spread,disseminated,
ifrån	off,
fiende	enemy,
grundlagen	constitution,the constitutional law,
odens	odin's,node,oden's,
universums	universe,the universe's,universe's,
pippi	birdie,pippi,
hamn	harbor,port,harbour,
nyare	newer,
knyta	tie,
kambodja	cambodians,
grönland	greenland,
status	status,
producera	produce,producing,
republikens	republic's,republic,
fysiologi	physiology,
protoner	protons,
persons	a person's,persons,person's,
linjerna	routes,the lines,lines,
göring	goring,cleaning,
producerad	produced,
vatikanstaten	vatican city,the vatican,vatican,
relaterade	related,
modet	the fashion,courage,fashion,
medvetna	aware,conscious,
kommunistisk	communistic,communist,
pennsylvania	pennsylvania,
breda	broad,qual o curso que você está estudando,wide,
hårdvara	hardware,hardwere,
without	without,
tjänsten	the service,service,
nordkoreas	north korea,north korea's,north coreas,
medellivslängd	average lifespan,life expectancy,
arkitekten	architect,the architect,
kopplingen	the connection,coupling,
lyckan	the happiness,happiness,
fördelas	be allocated,distribute,distributed,
listorna	menus,the lists of candidates,the lists,
kommentarer	comments,
förklarades	was explained,explained,
ekologiska	ecological,
enligt	according (to),according to,
kill	kill,
knäppupp	knäppup,knäppupp,
harrison	harrison,
märta	märta,
leta	search,check,
utvinns	extracted,
starka	strong,
tim	tim,h,
rose	rose,
regent	ruler,regent,
rosa	pink,rosa,
utbyte	yield,trade,
starkt	strongly,strong,
lett	resulted,led (to),
utvinna	extract,
pendeltåg	commuter train,commuter,
delstat	state,land,
feminism	feminism,
ross	ross,
riket	kingdom,the land,whole country,
mesta	most,
porto	postage,
vampyren	the vampire,vampire,
delhi	delhi,
utrikespolitik	foreign policy,foreign affairs,forgein policy,
uppslagsordet	lookup word,lexical entry; word,entry word,
kille	guy,
möts	meet,meets,
majoritet	majority,
inflation	inflation,
vampyrer	vampires,
walk	walk,
riken	the kingdoms,kingdoms,
kommentar	comment,
afrikas	africa's,africas,africa,
kennedy	kennedy,
höjer	rises,raise,raising,
cooper	cooper,
tower	tower,
anföll	attacked,
rammstein	rammstein,
verksamheten	the work,activity,
madrid	madrid,
innebära	mean,
teorin	theory,the theory,
gång	time,once,
passera	pass,
latinet	latin,
alkoholer	alcohols,
verksamheter	operations,businesses,activity,
försvarare	defenders,defender,
tiders	days',times,time's,
fiktion	fiction,
inspirerades	(was) inspired,inspired,
sitta	sit,
stopp	stop,
moon	moon,
härledas	derived,
lärda	literate,scholars,savants,
buddha	buddha,
lärde	learned,
uppbyggnad	construction,structure,
publicerat	published,
storhetstid	heyday,
liberala	liberal,
football	football,
servrar	servers,
geografi	geography,
genom	through,
tyskt	german,
korrekt	correct,
mandelas	mandelas,mandela's,
tyska	german,
tyske	german,
förbindelser	connections,relations,
on	on,
om	of,for,if,
indianska	red indian,amerindian,native american,
spelet	the game,game,
og	og,
of	of,av,
oc	o.c.,oc,
stand	stand,
hindu	hindu,
os	os,
spelen	the games,games,
befäl	command,
koppling	clutch,connection,
cambridge	cambridge,
ansträngningar	effort,
tolkning	interpretations,interpretation,
domstol	court,
överföras	transfer,transferred,
befinna	be,
mental	mental,
medlemsstaternas	member,member state,member states,
fisk	fish,
valley	valley,
serbien	serbia,
förrän	until,before,
genomfört	carried out,implemented,carried through,
flyga	fly,
inriktning	direction,orientation,alignment,
uppåt	raised,up,upwards,
ingredienser	ingredient,the ingredients,ingredients,
koenigsegg	koenigsegg,
manuskript	manuscript,script,
värre	worse,
ämbetsmän	officer,bailies,officers,
chaplin	chaplin,
kvinnornas	womens,the women's,women,
taylor	taylor,
felix	felix,
närmast	nearest,closest,mediately,
fjorton	fourteen,
pengar	money,
ökning	increase,
operation	operation,
köpenhamn	copenhagen,
många	many,
roses	roses,
mötley	mötley,
utgifter	expenditure,expenses,
babylon	babylonia,babylon,
visade	showed,showed; displayed,
separata	separate,
grupp	group,
sällskapet	society,the company,
symbol	symbol,
erövring	conquest,
missbruk	addiction,abuse,
vinnaren	winner,the winner,
observatörer	observers,
symtomen	symptoms,the symptoms,ymptoms,
villkor	conditions,condition,
distriktet	district,
barcelona	barcelona,
calle	calle,
erfarenhet	experience,
visby	visby,
all	any,
ali	ali,
alf	alf,
separat	seperate,separate,
samhället	the society,society,
stödde	supported,
samhällen	communities,societies,
utomliggande	external; ex-territorial,outlying,
sakrament	sacrament,
antogs	adoption,was assumed,
uppdrag	job,missions,mission,
persiska	persian,
funktionerna	functions,the functions,
brottet	offense,the crime,the crime; offense; infraction; transgression,
röstade	voted,
ögonen	eyes,the eyes,
gary	gary,
påstående	claim,assumption,
program	application,
cykeln	there are two meanings in the context - cycle and bicycle,cycle,
kvar	left,
löper	runs,at,
färgerna	colors,
woman	woman,
litet	small,
ansluter	connects,connect,
song	song,
far	father,
fas	phase,
fat	barrel,fat,
runtom	throughout,around,
simpsons	simpsons,
fan	devil,fan,
sony	sony,
redaktör	editor,
liten	small,
unionens	the union,european union,the union's,
tjeckiska	czech,
choklad	chocolate,
helvetet	hell,the hell,
list	cunning,
kopplas	connected,coupled,
förtryck	opression,
lisa	lisa,
programme	programme,
hitta	see,make up,come up, find,
grekland	greece,
ted	ted,
istiden	ice age,the ice age,
tex	for example,e.g.,
design	design,
haag	haag,the hague,
usama	osama,usama,
enklaste	the simplest,easiest,
sun	sun,
vaginalt	vaginal,
kinesiska	chinese,
version	version,
spelning	gig,playing,
sur	acidic,sour,
mördades	murdered,was murdered,murder was,
guns	guns,
fäste	bracket,attachment,
christian	christian,
dottern	the daughter,daughter,
upptäcka	detection,discover,
regerade	reigned,
avrättades	was executed,executed,
leeds	leeds,
madeleine	madeleine,
upptäckt	discovered,found,discovery,
norden	scandinavia; (nordic area; region),the nordic countries,north,
nordens	the scandinavian countries',scandinavia,nordic,
upptäcks	discoverd,detected,is discovered,
råder	advises,is,(that) prevails,
folktro	popular belief,folklore,
soloalbum	solo album,
kärnvapen	nuclear,nuclear weapons,
tillhörde	was a part of,belonging to,belonged to,
magnitud	magnitude,
arabemiraten	united arab emirates,uae,the arab emirate,
nyfödda	newborn,
påföljande	following,subsequent,
uppkomst	origin,onset,
kategorispelare	category player,
filmerna	films,the movies,
stöd	support,
syfte	purpose,view,
syfta	aim,refer,
smak	taste,flavoring,
socialdemokraterna	members of the social democracy,social democratic,
anarkism	anarchism,anarchy,
succé	succes,success,succession,
fängslade	inprisoned,confine,imprisoned,
branden	fire,the fire,
förebild	model,role model,
autonom	independent,autonomic,
bekräftade	confirmed,
genomsnittliga	average,
israel	israel,israeli,
permanenta	permanent,
cellerna	cells,the cells,
akademiens	academy,the academy's,attend,
glas	glass,
hålet	hole; gap,hole,the hole,
floyd	floyd,
glad	happy,
östra	eastern,
naturligt	natural,
legender	legends,
godkänt	approved,pass,
decenniet	decade,
gatorna	the streets,streets,
decennier	decades,
kryddor	spices,
förhåller	relate,relationship,relates,
naturliga	natural,
pony	pony,
division	division,
duett	duet,
bosatt	resident,lived,
huvudort	main town,principal town,
styrs	is controlled,ruled,
elektrisk	electric,elektirsk,
historiskt	historic,historically,historical,
court	court,
breaking	breakingpoint,breaking,
brittisk	british,
satanism	satanism,satanic,
historiska	historical,
härstamning	lineage,origin,descent,
välgörenhet	charity,
indelade	divided,divided into,
rocksångare	rock singers,rock singer,
skära	carve,cut,army,
sven	sven,
tagen	taken,
grundämne	elemental,element,
fötterna	feet,their feet,the feet,
ångest	anxiety,anguish,
fötts	born,borned,
atomer	atoms,
regnar	rains,raining,
anarkistiska	anarchistic,anarchist,
praktiska	practical,
bildade	formed,
tsar	tsar,czar,
homosexuella	homosexual,gay,
grande	grande,grand,
greklands	greece's,greek country,
människors	humans,human,people's,
friidrott	athletics,track and field,
längs	along,
avvisade	rejected,
september	september,
sträckte	extended,
emmanuel	emmanuel,
mission	mission,
australien	australian,australia,
längd	length,
retoriska	rhetorical,
hounds	hounds,
islam	islam,
lyder	reads,obeys,
rika	rich,
abbey	abbey,
rikt	target,rich,
prag	prague,
stephen	stephen,
argentina	argentina,
jämte	next (to),together with,plus,
fenomenet	the phenomenon,phenomenon,
kategorieuropeiska	european category,europe category,
styret	gate,
medborgerliga	civil,
kärna	core,quarks,
postumt	posthumous award,posthumously,
landborgen	the ridge,
marcus	marcus,
försöken	trials,attempts,the tries,
journalisten	journalist,the journalist,
krossa	crush,crushing,
stilen	style,
slidan	the vagina,vagina,vaginal,
journalister	journalists,
försöker	try,tries,trying,
principer	principals,principles,
kustlinje	coastline,
ringar	rings,
drycken	beverage,the drink,
betyg	grades,marks,
hawaii	hawaii,
konstnärlig	art,artistic,
aldrig	never,
drycker	beverages,
stenar	stones,blocks,
ollonet	penis head,glans,the glans,
därvid	thus; thusly; then,therewith,in so doing,
nepal	nepal,
europas	europe,
hill	hill,
väg	vague,way,
kvinna	woman,
väl	selecting,good,
vän	van,friend,
benjamin	benjamin,
poliser	police (-men; -women),police,
ökad	increase,increased,
islamistiska	islamic,islamist,
densiteten	density,
beräknades	calculated,estimated,
kritiserat	criticized,criticised,
spelades	filmed,
kritiserar	criticize,
polisen	police,the police,
faller	fall,
fallet	case,the case,
stavningen	spelling,the spelling,
konsumtionen	the consumtion,consumption,
fallen	case,cases,
aminosyror	amino acids,
filosofins	philosophy,the philosophy,
heinz	heinz,
colombia	colombia,
pablo	pablo,
bland	blamd,inter,including,
blanc	blanc,
story	story,
infört	introduced,
lördagen	the saturday,saturday,
automobile	automobile,
misslyckas	fail,fails,
harris	harris,
stort	large,big,
motiveringen	the motivation,ground,
storm	storm,
kristendomens	christianity's,the christianity's,christianity,
brasiliens	brazil's,
ecuador	ecuador,
familjerna	families,
mikael	mikael,
gränser	borders,frontiers,
hotel	hotel,
kongress	congress,
serotonin	serotonin,
framtiden	future,the future,
hotet	the threath,the threat,threat,
fattigaste	the poorest,poorest,
gränsen	limit,border,the line,
besökare	visitors,
siffra	number,figure,
king	king,
illegala	illegal,irregular,
matcherna	the games,games,
direkt	direct,directly,
kina	china,
pjäsen	play,piece,
dans	dance,
kategorisommarvärdar	category summer hosts,
guden	god,the god,
stjärnan	star,the star,
tillåta	allowing,allow,
klubb	club,
anläggningar	plants,facilities,
kusin	cousin,
tilldelas	assigned,award,
tabell	table,chart,tabel,
omskärelse	circumcision,
slåss	fight,
divisionen	division,
wilson	wilson,
bakgrunden	background,
bedriver	conducts,manage,operate,
inriktningar	direction,specializations,
dialekt	dialect,brogue,
jämförelsevis	comparative,in comparison,comparatively,
judas	judas,
judar	jews,
kiss	kiss,view,
folkgrupper	communities,ethnic groups,
electric	electic,electric,
dagliga	daily,
park	park,
stjärnans	star's,the star's,the stars,
dagligt	daily,
industrialiserade	industrialized,
agnostiker	agnostic,agnostics,
sånger	songs,
mineral	minerals,mineral,
windows	windows,
salt	salt,
influensan	the influenza,flu,
sången	the song,song,
zeppelin	zeppelin,
statsskick	polity,form of government,government,
kosovo	kosovo,
tjugo	twenty,
rösta	vote,
ursprungliga	original,
kapitulerade	surrendered,
tilly	tilly,
månen	the moon,man,
förening	union,compound,
beräkningar	calculations,
canaria	canaria,
grace	grace,
moses	moses,
his	his,
hit	to here,here,
hiv	hiv,
stormakterna	great powers,
inklusive	including,
vardera	either,each,
b	b,
jobbade	worked,
händer	happens,happening,hands,
sofie	sofie,
solsystemet	the solar system,solar system`,
budapest	budapest,
utvidgade	expanded,
tvkanaler	tv-channels,tv channels,
mediciner	medicines,
avtal	agreement; deal,agreement,contract,
tidszon	timezone,time zone,
vincent	vincent,
norrköping	norrköping,
poäng	score,point,
virginia	virginia,
utsatt	exposed,
bars	bar,carried,
etiopien	ethiopia,ethiopian,
art	kind,art,
bart	offense,bart,
arv	heritage,
fiske	fishing,
bara	only,
are	are,
arg	angry,
flyttade	moved,
stjäla	steal,stealing,
arm	arm,
barn	child,
pär	pär,
bortsett	except,apart,
planeras	is planned,planned,
överföring	transfer,
uppskatta	estimate,appreciate,
inga	not,no,
planerat	planned,
invaldes	elected,was elected,
planerad	planned,
oerhörd	tremendous,
verksamhet	work,activity,
där	where,in which,were,
intäkter	revenues,incomes,
herrar	gentlemen,men,
uppkom	arose,
godkändes	was approved,approved,
tiderna	the times,times, ages,time,
balkanhalvön	balkans,balkan peninsula,
startades	started,
operan	opera,the opera,
roman	novel,
lägret	the camp,camp,
påstår	states,claims,asserts,
hypotesen	the hypothesis,hypothesis,
lära	lara,get to know,learn,
borta	gone,away,
vidare	moreover,furthermore,further,
lärt	learned,learnt,
stärktes	was strengthened,strengthened,was strenghten,
belägna	located,disposed,
besegrade	defeated,
östtyskland	east germany,
utifrån	from the outside,from,
hypoteser	hypotheses,hypothesis,
ps	ps,p.s,p.s.,
java	java,
göteborg	gothenburg,
personalen	personnel,the staff,
kungafamiljen	the royal family,
johannes	johannes,john,
avslutade	ended,finished,
byxor	pants,
resultat	results,result,
ph	ph,
pi	pi,
chandler	chandler,
flight	flights,flight,
togs	taken,were taken,
publiken	the audience,audience,
sydafrikas	of south africa,south african,south africa's,
rättigheterna	the rights,rights,
gården	farm,courtyard; house; farm (-house),
konflikter	conflicts,conflict,
konflikten	the conflict,conflict,
deltog	participated,
julius	julius,
sådan	such,kind of,
inspelningar	recordings,
ägs	is owned,(is) owned,owned,
styr	controls,
ris	rice,
rik	rish,rich,
sjöarna	the lakes,lakes,
byggnaderna	building,buildings,the buildings,
skeppen	the ships,
fysisk	natural,physical,
demografi	demographics,demography,
tidpunkten	the time,the moment,time,
ideologier	ideologies,
sjunkit	decreased,
förföljelse	persecution,
torbjörn	torbjörn,torbjorn,
spears	spears,
låtit	had,let,ordered,
bröllopet	the wedding,wedding,
byar	villages,
skåne	skåne,scania,
uppbyggd	structered,structured,built-up,
författare	author,
uppbyggt	structured,
kokpunkt	having a boiling point,boiling point,
vinklar	angle,angles,
finansiera	fund,finance,
italiensk	italian,
sjunga	access,sing,
edge	edge,
vetenskapen	the science,science,
kyrkans	the church's,the churche's,church,
alfabet	alphabets,alphabet,
uttalande	statement,
kontinentala	continental,
komplett	complete,
konstitution	constitution,
påverkade	influenced,affected,
remmer	remmer,
dåtidens	past times,yesterdays,that time,
prince	prince,
namnet	name,the name,
folkräkning	census,head count,
skalv	shock,quake,
minoriteter	minorities,
bostad	lodge,property,
omedelbar	instant,immediate,
försvunnit	disappeared,
skall	is,shall,
centralasien	central asia,
idé	regard,ide,
emigrerade	emigrated,
px|centrerad	px | centric,
skala	scale,scale; size,
färdiga	finished,completed,
synnerhet	specially,particular,
djupare	depth,deeper,
rastafarianerna	the rastafarian,rest are faria,n/a,
begravdes	buried,
användas	used,
stoppade	stop,stopped,
upplevelse	experience,
exakt	precise,accurately,
våldsamma	violent,
näringsliv	business,
banbrytande	groundbreaking,
sammansättning	composition,
hittar	found,finds,
hittas	found,be found,
hittat	found,
minskning	decline,reduction,decrease,
landskommun	rural municipality,
norrut	north,
sjöfart	sea voyage,navigation,maritime,
kongo	congo,kongo,
lettland	latvia,
trummis	drummer,
global	global,
krigare	warriors,warrior,
flottan	the fleet,navy,the navy,
thailand	thailand,
huvudstad	capital city,capital,
låtarna	the songs,songs,
ungefär	approx.; approximately,about,approximately,
höjden	height,
föräldrar	parents,
grekerna	greeks,greek,
prov	test,tests,
frälsning	salvation,
fungera	act,
anne	anne,
trinidad	trinidad,
höjdes	increased,was raised,
höjder	altitudes,heights,
turism	tourism,
diamant	diamond,
palmes	palme,palme's,plame's,
ställningen	position,
tävlade	competed,
presenteras	was presented,presented,
anklagades	accused,
bayern	bavaria,bayern,
judendom	judaism,jewism,
kostnaderna	costs,the costs,
grundläggande	because lag of,primary,fundamental,
påtryckningar	pressure,pressures,
tätt	tight,tightly,
virus	virus,
ande	of,spirit,
dialog	dialogue,
täta	close,seal,
socialistisk	socialistic,socialist,
oktoberrevolutionen	the october revolution,october revolution,
genomföras	carried out,be performed,carry out,
medborgarna	the citizens,citizens,
reglerna	rules,rules; regulations,
hållet	cohesive,way,
abbas	abbas,
km²	square kilometre,km2,
laget	the team,stroke,
håller	is,holds,
dricka	drinking,drink,
long	longitude,long,
jugoslavien	yugoslavia,
bagge	bagge,ram,
bruk	using,use,
laila	laila,
ateister	atheists,steister,
delning	division,pitch,
rasade	collapsed,
regionen	the region,region,
längtan	longing,
sköter	handles,handle,
kritikerna	critics,the critics,critiques,
delta	participate,delta,
regioner	regions,
junior	junior,
medeltidens	ages,medieval,
anklagelser	allegations,accusations,
planeternas	the planets,planets,the planets',
världskrigen	the world wars,world wars,
styrande	rulers,governing,
aktier	share,stock,
erövrades	conquered,(was) conquered,concoured,
guyana	guyana (name),guyana,
tolka	interpreting,interpret,
handels	commercial,trade,
z	z,
tidens	time's,time,that time's,
svenskspråkiga	swedish speaking,swedish-speaking,
ägdes	owned,
singlarna	singles,the singles,
tidpunkt	date,time,
home	home,
däribland	among them,including,
graham	graham,
veckorna	weeks,
rainbow	rainbow,
stadion	stadium,the stadium,
möten	meetings,
höga	high,
psykoterapi	psychotherapy,treatment,
högst	highest,maximum,
mötet	the meeting,meeting,
hanen	the cock,the male,male,
urval	selection,
skyddas	protected,(is/are) protected,
skyddar	protection,protects,
sutra	sutra,
beräknas	calculated,estimated,
beräknar	calculates the,computes,values,
tittarna	the viewers,viewers,
medina	medina,
stadigt	stable,steadily,
konvertera	conversion,convert,
betyder	means,
råkar	happens,happens to,
kaspiska	caspian,
modernismen	modernism,
klubbens	club,
oväntat	unexpectedly,unexpected,
underlättar	make it easier,facilitates,
vice	vice,
europeiska	european,
parallella	parallel,
microsoft	microsoft,
nasa	nasa,
karma	karma,
lagstiftning	law-making,regulation,
europeiskt	european,
nash	' nash,nash,
förhandla	negotiate,negotiating,
psykologi	psychology,
beträffande	on,
kanal	channel,
steve	steve,
jimi	jimi,
stieg	stieg,
moseboken	genesis,
norrköpings	norrköpings,
simon	simon,
uppmaning	call; injunction,call,exhortation,
fortfarande	still,
romerna	the romani people,the romani,roma,
kazakstan	kazakstan,kazakhstan,
generellt	generally,
generella	overall,general,
hinduism	hinduism,
fotnoter	footnotes,
pengarna	the money,money,
varierar	varies,vary,
vapen	weapons,weapon,
kategoritvseriestarter	category television series starts,
varierat	varied,
mesopotamien	mesopotamia,
sjukdomar	diseases,disease,
medverkade	participated; contributed,participated,
kommitté	committee,
avslutas	close,ends,closing,
avslutat	completed,finished,
tvinga	force,
historikern	historian,the historian,
paz	paz,
demokratiskt	democratic,
markera	mark,
inleder	start,initiates,
noter	notes,notation,
byggs	building,under construction,
sällsynt	rare,
utanför	outside,
melodier	melodies,
byggd	built,
demokratiska	democratic,
bygga	building,build,
indirekt	indirect,indirectly,
skadad	damaged,
åtminstone	at least,
århundradet	century,
skadan	damage,the damage,the hit,
influerad	influenced,
anderssons	anderssons,andersson's,
skadas	damaged,
västlig	western,
konstant	constant,
folk	public,people,
influerat	influenced,
hölls	was held,was,
assisterande	assistant,assisted,assisting,
kris	crisis,
skrivna	written,
domkyrka	cathedral,abbey,
krig	war,
dramatiska	dramatic,dramatical,
bröts	was fractured,broke,
koloni	colony,
hdmi	hdmi,
producenten	the producer,producer,
turismen	tourism,the tourism,
producenter	producers,
diamanter	diamonds,
åtgärder	measures,
filosofi	philosophy,
astrid	astrid,
tvingats	forced,had,
fauna	fauna,
buddhistiska	buddhistic,buddhist,
ukraina	ukraine,
metro	metro,
innehar	holds,holding,
innehas	held,occupied,
innehav	possession,holdings,owning,
springsteens	springsteen's,springsteens,
plattan	plate,the plate,
fortsätter	continues,continue,
populärkulturen	popular culture,
översättningar	translations,
tjänar	earns,serves,
zlatan	zlatan,
reda	find out,out,find our,
gemenskap	fellowship,community,
föreställande	depicting,
motor	engine,
juryns	the jury's,jury,
redo	ready,prepared,
varpå	thereafter,whereupon,after which,
from	from,
bestämmelser	regulations,measures,conditions,
usa	the usa,united states of america,usa,
fel	faults,errors,error,
fem	five,
sevärdheter	attractions,
upplöstes	dissolved,
källorna	source,the sources,
inlandet	inland,the inland,
öppnat	opened,opening,
andliga	spiritual,
penis	penis,
införande	introduction,
hindrade	preventing,prevented,
vägrade	refused,
fungerar	functions,works,
reguljära	regular,
beskriva	describe,
automatiskt	automatic,
beskrivs	described,
tar	takes,
tas	is,is taken,
föreslår	suggests,suggest,
ledamöterna	the commissioners,commisioners,the members,
crick	cricket,crick,
engels	engels,
treenigheten	tinity,the trinity,trinity,
tag	while,
hilton	hilton,
tal	speech,
kanadensiska	canadian,
sir	sir,
omvänt	reversed,vice versa,
löften	promises,
beyoncé	beyonce,beyoncé,beyoncè,
six	six,
brian	brian,
sig	to,itself,
undantaget	except,
sin	its,
väpnad	armed,
kostym	costume,
kontroversiellt	controversial,
förekommande	occuring,where,
oavsett	whether,regardless; whether; irrespective of,regardless,
tack	thanks,
religiös	religious,
bertil	bertil,
kategoriwikipediabasartiklar	category wikipedia basartiklar,
kontroversiella	controversial,
eritrea	eritrea,
light	light,
centralorter	centers,regional centers,
framförts	forward,performed,
öresund	Øresund,the sound,
jolie	jolie,jolies,
besegrat	defeated,
mekka	mecca,mecka,
blandad	mixed,blended,
skapande	building,creating,creative,
företrädare	representatives,
elin	elin,electrical,
förklaras	explained,
elit	elite,
blandat	mixed,
karlstad	karlstad,phoenix,
blandas	mixed,mixes,
spotify	spotify,
stiga	rise,rising,
uppmärksammad	noted, come to attention,attention,noticed,
terriers	terriers,
befolkning	population,
byn	village,
floder	rivers,
permanent	permanent,
försvar	defence,defense,
datorn	the computer,pc,
thåström	thåström,thastrom,
carola	carola,
skede	period,analysis,
cypern	cyprus,
verkligen	real,the reality,
washington	washington,
fler	more,
östtimor	east timor,
satelliter	satellite,
exempelvis	e.g.,
komma	access,get,
ale	ale,
billy	billy,
växande	growing,
konungariket	kingdom,
vidta	take,
studios	studios,the studio's,
boende	resident,housing,accommodation,
säsonger	seasons,
barnets	the childs,the child's,child,
byter	changing,changes,exchanges,
kvarteret	quarter,the neighborhood,
säsongen	season,
studion	studio,the studio,
kritik	criticism,critisism,critique; criticism,
alger	algaes,algae,
förbjuda	forbid,ban,prohibiting,
uggla	owl,
minskad	decreased,reduced,
hantverkare	handy worker,craftsman,
fiktiva	fictitious,romantic,
svar	answer,response,
bål	prom,torso,
nobelpristagare	nobel laureate (-s); nobel prize winner (-s),nobel laureates,
minskat	decreased,reduced,has decreased,
uppnå	achieving,achieve,
minskar	diminishing,decrease,
förutsättningar	prerequisites,(pre-)conditions,condition,
hörs	heard,
hört	heard,heared,
hjälpt	helped,
vulkanutbrott	vulcano eruption,volcanic eruption,
utmärker	characterizes,characterized,
höra	hear,know,
hjälpa	helping,
york	york,
studioalbumet	studio album,
philip	philip,
domare	judge,
hörn	corner,
fotbollslandslag	football team,national football team,
gångna	past,past; gone,
anslutning	connection,
tyst	quiet,silent,
waterloo	waterlo,waterloo,
g	(g),
barns	child,childrens,children,
via	via,through,
adrian	adrian,
tvserier	tv-shows,tv shows,tv-series,
tysk	german,
rudolf	rudolph,rudolf,
ovanpå	top,on top of,
revolutionens	revolution,the revolutions,
isbn	isbn,
brasilien	brazil,
velat	wanted,
kriterier	criteria,
värsta	worst,
mått	measurements,measurement,measure,
skyddade	protected,
nätverk	network,
enkelt	simple,easy,
förhöjd	enhanced,elevated,
fågelhundar	bird dogs,
meddelanden	messages,
omfattning	extent,
misslyckande	failure,
sankta	sankta,saint,
diskutera	discussed,discuss,
rösträtt	vote,right to vote,
valde	crowned,selected,chose,
valda	chosen,
vingar	wings,
juli	july,
vind	wind,
dödligheten	mortality,
institution	institution,
franska	french,
holland	holland,
franske	the french,french,
birgitta	birgitta,
tommy	tommy,
framgång	success,
algeriet	algeria,
franskt	french,
tomma	empty,
tyskarna	the germans,germans,the german,
distinkt	distinct,distinctive,
fyrtio	forty,
cohen	cohen - it's a name,cohen,
benny	benny,
avgörs	determined,is determined,decided,
blir	become,is,
farligt	dangerous,hazardly,
ringen	ring,
gäng	group,thread,
intervju	interview,
storbritannien	great britain,uk,
byggas	prevented,built,build,
uppfann	invented,
lopp	course, passage,races,race,
ansåg	thought,found,considered,
besittning	dominion,possess,
kristi	kristi,christ,
betydligt	considerably,significant,
centra	center,
ström	stream,power,icon,
centre	center,centre,
who	who,
intogs	was taken,was captured,
representation	representation,
staternas	states,the state's,
öken	desert,
planerade	planned,
förbundsrepubliken	the federal republic,federal republic of,federal republic,
undersökte	investigated,examined,
regeringschef	head of government,government,
miljontals	millions,
enbart	only,
judendomen	the judaism,judaism,
kategoriamerikanska	u.s. category,
movie	movie,
moberg	moberg,
uefa	uefa,
blandade	mixed,
funktionella	functional,
debatt	debate,
julafton	chistmas eve,christmas eve,
pastoral	pastoral,
angående	concerning,reference,
dödades	killed,were killed,
asterix	asterix,
rösten	voice,rust,the voice,
filmer	films,movies,
röster	votes,
beroende	dependent,dependent on,depending,
hållning	position,attitude,entertainment,
allmänhet	in general,public,general,
träffa	meet,see,
gränsar	border,adjacent,borders (to),
heta	hot,be named; be called,be called,
samtida	contemporary,
gudar	gods,
linje	line,
presley	presley,
hett	hot,
närstående	relative,relatives,kindred,
samtycke	consent,approval,
städer	urban,cities,
begäran	request,
förbinder	connects,undertake,
torka	dry,
respektive	and,respective,
mestadels	most of the time,mostly,
kvinnorna	the women,women,
berömd	famous,
nationernas	the nation's,the nations,nations,
rikare	richer,
motståndare	opponents,opponent,
ansågs	was,seemed,
funktion	function,
upplysning	the enlightenment,enlightenment,
praktisk	practical,
sydstaterna	the southern states,southern states,southern united states,
faktiskt	in fact; actually; indeed,really,actually,
vandrar	wanders,migrates,
joe	joe,
swift	swift,
jon	jon,
sångaren	singer,the singer,
allsvenskan	headlines,allsvenskan,
ingemar	ingemar,
påtagligt	substantially,considerably,markedly,
utvecklingen	development,the development,
teoretiker	say,theorists,
kolhydrater	carbons,carbohydrates,
april	april,
västerländsk	western,
brons	bronze,
vattnets	water,the water's,the waters,
bronx	bronx,the bronx,
klasser	classes,
betecknar	represent,denotes,represents,
betecknas	designate,labelled,denote,
kategorityska	category: german,
exakta	exact,
korruption	corruption,
wall	wall,
vittne	witness,
publicerad	published,
walt	walt,
cirka	about,approximately,
utsedd	appointed,
styrkor	strenghts,forces,
publiceras	publishes,will be published,published,
framträdanden	appearances,
jenny	jenny,
utkom	issued,(was) issued,published,
klara	clear,
dödshjälp	euthanasy,euthanasia,
nåddes	reached,
kopplade	connected,
bbc	bbc,
beskrivning	description,
månar	moons,
marilyn	marilyn,
klart	clear,done,finished,
månad	month,
strindbergs	strindberg's,strindberg,
ständig	constant,
naturtillgångar	natural resources,
mike	micke,mike,
liverpool	liverpool,
nickel	nickel,
klassen	the class,
turneringen	the tournament,
dominera	dominate,
lutherska	lutheran,
försvann	disappeared,
hms	hms,
fortsättningen	the continuation,remain,
neutrala	neutral,
deklarerade	declared,
last	load,
plikter	duties,
present	gift,
godkännande	approval,authorization,
bråk	brawl; fight,fights,fraction,
problemen	problems,the problems,
officiell	official,authentic,
största	biggest,maximum,largest,
anpassa	adjust,adapt,
will	will,
fördelade	divided,distributed,
yngre	younger,
wild	wild,
fjärdedel	quarter,fourth,
värmlands	varmlands,värmlands,hot countries,
explosionen	the explosion,
sagan	story,
uppfattning	understanding,view,
gemensamt	single,in common,
bosättare	settlers,
syftar	refers,seek to,refer,
motiv	subjects,motif,
jehovas	jehovas,jehova's,
röra	move,
uppstå	develop,occur,arise,
ramels	ramel's,
varar	duration,lasts,
buddhism	buddhism,
pojkar	boys,
samband	connection,
inch	inches,
skickade	sent,
gett	given,gave,
annekterade	annexed,annexation,
tvister	conflicts,disputes,
mottagande	host,reception,
övervägande	the predominant,predominant,predominantly,
romeo	romeo,
romer	romani people,roma,
student	student,
raka	straight,
rätt	right,entitled,
misstag	error,mistake,
klubbar	clubs,
vilar	rests,
banden	bands,bander,the bound,
terrorismen	terrorism,the terrorism,
undersökningar	surveys; investigations,studies,studies',
närma	approach,move closer,approximate,
ekosystem	ecosystem,eco system,
övertyga	convince,
english	english,
bandet	band,
organisationens	organization,the organizations,
hårdrocken	hard rock,
lön	salary,wage; salary,
biologisk	biological,
singeln	single,singeln,
mfl	etc,etc.,
möjligheter	potential,
uppkommer	arises,resulting,arises; generated,
möjligheten	the ability,the possibility,
rachels	rachels,rachel's,
erfarenheter	experiences,experience,
högskolor	colleges,
patrik	patrik,
miljöer	environment,environments,
antisemitism	antisemitism,
rocken	the rock,rock,
brutit	cut; break,broken,
mytologiska	mytholigical,mythological,
jarl	earl,jarl,
genombrottet	break-through,breakthrough,
alldeles	completely,altogether,
hoppa	skip,drop out,
bell	bell,
sky	sky,
rättsliga	justice,legal,
engelsk	english,
ske	be,happen,
ska	will,shall,
fyller	turns,play,turn; fill,
sanskrit	sanskrit,
hotade	threatened,
psykoser	psychoses,psychosis,
färgen	color,the color,
olle	olle,
agerande	acting,behavior,
älska	love,
know	know,
press	press,
psykosen	psychosis,the psychosis,
säljs	sold,
georges	georges,
budet	the bid,the commandment,
miami	miami,
djupa	deep,
huruvida	whether,
sälja	sell,
gorbatjov	gorbachev,gotbatjov,
immunförsvar	immune,immune defense,
finansieras	financed,funded,finansed,
djupt	deeply,deep,
säkra	reliable,safe,secure,
serbiska	serbian,
tjeckoslovakien	czechoslovakia,
handeln	trade; commerce,trade,
berömt	famous,praised,
bibliska	biblican,biblical,
efterfrågan	demand,
gäst	guest,
export	export,
försvinna	vanish,disappear,
star	star,
empire	empire,
skandinavien	scandinavia,
använts	was used,used,
genomsnitt	average,
planering	planning,
trianglar	with triangles,traingles,
gammalt	old,
tvfilm	tv-movie,tv film,tv movie,
undviker	avoids,avoid,
klassificera	classifying,classify,
setts	observed,seen,
mankell	mankell,
låter	let,
låten	the song,song,
sjunker	flag,sinks,
äta	eat,
utsöndras	secrete,exudes,secreted,
uppvärmning	heating,warming,
mitt	my,center,
slut	end,out,
dateras	dates,dated,
sommarspelen	summer games,summer olympics,
lång	long,
ljung	heather,
låna	borrow,lana,
koalition	coalition,
substantiv	noun,
tillräcklig	sufficient,enough,
överlevde	survived,
bestämma	determining,decide,
oberoende	independent,
avsnittet	section,episode,
saken	the thing,matter,the matter,
saker	things,items,
avsnitten	the episodes,sections,chapters,
mäta	compare,feeding,
own	egen,
främre	forward,front,
egna	own,custom,
återvänt	returned,returning,
någorlunda	fairly,somewhat,
avrättade	executed,
tillbringade	spent,
mäts	measured,is measured,
sektorn	sector,the sector,
floden	river,the river,
mätt	measured,dull,
flyger	flies,flying,
stressorer	stressors,
glukos	glucose,
folkpartiet	peoples party,liberal party,
konstruktion	construction,structure,
födelsetal	birthrate,birth rate,
citat	quote,
val	choice,elections,election,
idén	the idea,idea,
vad	as,what,
smeknamnet	nickname,
mäter	measuring,measure,
var	was,
regisserad	directed,produced,
bevarade	preserved,
nordamerikanska	north american,
lundell	lundell,
granne	neighbour,neighbor,
hundratal	100,hundred,
ingått	been part of,entered,entered into,
krigsslutet	end of war; war's end,end of the war,
stadens	the town's,the citys,city's,
karta	map,maps,
made	made,
rybak	rybak,
arne	arne,
tema	theme,
missnöjet	discontent,grievance,
kuriosa	bric-a-brac,curiosities,trivia,
reaktorn	the reactor,reactor,
problemet	problem,the problem,
stormakter	world powers,great power,superpowers,
eu	eu,
utöva	carry,utÖva,exercise,
runor	runes,
kant	kant,edge,
året	the year,all year,years,
illinois	illinois,
rike	kingdom,
book	book,
ursprunget	origin,the origin,
åren	the years,years,
intresse	interest,
juni	june,
tillhörighet	affiliation,belonging,belonging; affiliation,
tolkas	is interpreted,interpretation,interpret,
tolkar	interprets,views,
shakespeares	shakespeare's,shakespeare,
risker	risk,risker,risks,
personligen	individual,personally,
taube	taube,
ställningar	positions,standings,notions,
margaret	margaret,
markant	considerably,markedly,marked,
risken	the risk,risk,
cliff	cliff,
nödvändigtvis	by necessity,necessarily,
knappast	hardly,dead,
inledning	introduction,the beginning,
bysantinska	byzantine,
blogg	blog,
tidning	newspaper,journal,
