vanligast	most usual,
nordisk	norse,nordic,
uppemot	almost,
stammarna	tribes,
arternas	the species,
jihad	johad,jihad,
elva	eleven,
invandrare	immigrants,
hållas	be held,
albumet	album,
slå	hit,
albumen	the albums,
hermann	hermann,
lord	lord,
vann	won,
lyckats	succeeded,
dela	divide,
syrgas	oxygen,
regional	regional,
upptar	occupies,
lämnades	left,
portugals	portugal,
dels	both,
skicklig	skillful,skilled; skillful,
statlig	government,
medelhavet	mediterranean sea,
andre	other,
helsingborg	helsingborg,
haber	haber,
befogenheter	authorities,
triangelns	the triangle's,
urskilja	distinguish,discern,
sovjetisk	soviet,sovjetic,sovietic,
miller	miller,
sture	sture,
sammansatta	composite,composed,joined,
selassie	selassie,
ungerns	hungrarys,hungary's,
hanar	males,
upprätthåller	maintains,
åsikten	the opinion,
åsikter	opinions,
breddgraden	latitude,
fossil	fossil,
punkt	point,
jönsson	jönsson,
filosofer	philosophers,philosopher,
aten	athens,
hårda	hard,
biografi	biography,
vägrar	refuses,refuse,
filosofen	the philosopher,
motståndsrörelsen	the resistance,resistance,
regnskog	rain forest,
analytisk	analytical,
föräldrarna	the parents,
valrörelsen	election campaign,
bipolär	bipolar,
kids	kids,
demokratier	democracies,
naturen	the nature,nature,
blåser	blows,blowing,
vicepresident	vice president,
robin	robin,
miljarder	billions,
systematiska	systematical,
unik	unique,
norsk	norwegian,
välkänd	well-known,well known,
hamas	hamas,
systematiskt	systematically,systematic,
ansluta	join,connect,
dna	dna,
sjukdomen	disease,
strikt	strict,
fuktiga	damply,
betraktats	considered,been seen,(been) viewed,
 mm	millimeter,
dns	dns,
fuktigt	moist,humid,
musik	music,
dickens	dicken's,
befolkningstillväxten	population growth,the population growth,the growth of population,
mercurys	mercury's,mercurys,
holm	holm,
politiker	politician,
slutligen	finally,
bulgariska	bulgarian,
kalksten	limestone,
teman	themes,
ofta	often,
vännen	the friend,friend,
köpa	purchase,buy,
befolkningsutveckling	population development,
vågen	the wave,
stommen	frame,the foundation,
köpt	purchased,bought,
passagerare	passenger,
kapitalismen	capitalism,
want	want,
absoluta	absolute,
vänner	friendas,friends,
hon	she,
kallare	colder,
hov	court,
how	how,
pågick	lasted,
folkmusik	folk music,
typen	model,the type,type,
fylla	fill,
inrikes	domestic,
trettioåriga	13 year olds,thirty year's (war),
barbro	barbro,
sedd	seen,
objekt	objects,
turkiet	turkey,
sankt	st.,sankt,
typer	characters,types,
stormaktstiden	great power period,
grekiska	greek,
isär	apart,
arbeten	works,
hemlandet	the homeland,
wind	wind,
skådespelerska	actress,
varv	dockyard,shipbuilding,
dahléns	dahlén's,
vars	who's,
dalí	dali,
organismen	the organism,
vare	either,
varg	wolf,
organismer	organism,
vara	be,
barnet	child,
mabel	mabel,
varm	warm,
publicerade	published,
besläktade	related,
nutida	present(-day); contemporary,present day,
wales	wales,
assyriska	assyrian,
avgå	resign,
väte	hydrogen,
säljande	selling,
bestämmer	determines,decide,
hänga	hang,
närliggande	nearby,
silver	silver,
utvecklat	evolved,
utlänningar	foreigners,
utvecklar	develops,
framsteg	progress,
terrorister	terrorists,
tingslag	leet,
debut	debut,
utveckling	development,
tillgängligt	available,
utvecklad	developed,
tillgängliga	available,
uppnådde	achieved,
talade	spoken,
lätt	easy,
serier	comics,
allan	allan,
kontroverser	controversies,contraversies,
serien	series,the series,
avståndet	the distance,
axelmakterna	the axis,axis,
varken	neither,either,
kontrollerade	controlled,
försökt	tried,
förändringar	changes,
snarare	rather,
anarkister	anarchists,
metallica	metallica,
arbetsplats	work,workplace,
ägnade	dedicated,
sannolikt	probable,
att	to,that,
sysselsätter	employs,
okända	unknown,
malmös	malmö's,
sydost	south east,
givetvis	naturally,
grannlandet	the neighbouring country,
östberg	Östberg,
tecknade	cartoon (-s),cartoon,drew,
övre	upper,
ledarskap	leadership,
förespråkar	advocate,
xis	the eleventh's,
master	master,
vågade	dared,
ära	glory,
bitter	bitter,
förändringarna	changes,
senaten	senate,the senate,
bokstäverna	the letters,
förmögenhet	wealth,
placerade	put,placed,placed (in),
leukemi	leukemia,
nirvana	nirvana,
påverkad	influenced,affected,
ahmed	ahmed,
skatter	taxes,
upphov	origin,source,
tyckte	thought,
påverkan	impact,influence,
tree	tree,
upplysningstiden	enlightenment,age of enlightenment,
nations	nations,
trey	trey,
varje	each,
utformningen	the layout,layout,the design,
påverkas	affected,
tretton	thirteen,
obligatorisk	obligatory,mandatory,
försörja	support,
boston	boston,
dricker	drink,drinks,
filosofisk	philosophic,
albanska	albanian,
joakim	joakim,
trakten	the region,region,
fasta	firm; set; solid; fast; fasting,
kroatien	croatia,
normalt	normally,normal,
östeuropa	eastern europe,east europe,
skaffa	get,
förhärskande	dominant,prevailing,
himlen	heaven,although the sky,
hjälpmedel	aid,resources,
bedrivs	conducted,
katalonien	catalonia,
konserthus	concert hall,
victoria	victoria,
gallagher	gallagher,
medlemsstaterna	member states,
anteckningar	notes,
bedriva	prosecute,
eftersom	while,because,
thriller	thriller,
övertog	took over,overtook,
singer	singer,
morgon	morning,
arkitektur	architecture,
hämnd	revenge,
camp	camp,
utmärkande	distinguishing,
förlorar	loses,
översatt	translated,the translation,
förlorat	lost,
konstantinopel	constantinople,
passerade	passed,
singel	single,
tänkte	thought,was going to,
majs	corn,
ungar	babies,kids; offsprings; young,
representanter	represenatives,representatives,
bomb	bomb,
bandmedlemmar	band members,
diplomatiska	diplomatic,
nacka	nacka,
legitimitet	legitimacy,
teater	theatre; theater,theater,
louise	louise,
populärkultur	popular culture,pop-culture,
buss	bus,
övergår	surpasses,released,exceed,
sekulär	secular,
bush	bush,
omvända	reverse,
mottog	received,
lastbilar	truck,trucks,
tillståndet	condition,the state,
rättegången	the trial,
årsdag	anniversary,
metoder	methods,
upprätta	establish,
metoden	the method,
dansk	danish,
plats	place,spot,place; position,
nathan	nathan,
lyssna	listen,
begravning	funeral,
hantverk	crafting,
×	x,
kallt	cold,coldly,
sköta	manage,operate,handle,
roy	roy,
utgåvan	edition,issue,the edition,
uppgift	task,
genomsnittet	average,the average,
sköts	postponed; run,handled,
kalla	cold,
blev	became,
etik	ethics,
flagga	flag,
skulle	could,would,
skriva	write,
bygger	(is) building (on),
arlanda	arlanda,
skrivs	written,
nuförtiden	today,
hedersdoktor	honorary doctor,honorary degree,
manson	manson,
förhindra	prevent,
wikipedia	wikipedia,
upphovsrätt	copyright,
sundsvalls	(city of) sundsvall's,
sista	last,
siste	last,
österrike	austria,
ringa	call,
rollen	the role,
henrik	henrik,
ställning	position,
lanserades	launched,
konsekvens	consequence,
tilldelades	awarded,
kommunikation	communication,
världsturné	world tour,
roller	roles,
tillämpar	administer,practice,administers,
huvudet	head,the head,
kubas	cuba's,
följas	followed,
pitt	pitt,
nordiska	nordic,
nederlag	defeat,
nordiskt	nordic,
genus	genus,
logik	logic,
aktuell	current,
igelkotten	the hedgehog,hedgehog,
folkmordet	genocide,
armén	the army,
uttal	pronunciation,
herr	mister,mr,
ana	feel,
union	union,
avgörande	settling,decisive,
fri	free,
anc	anc,
operationer	operations,
socialistiskt	socialistic,socialist,
årtionde	decade,
fru	madam,wife,
arbetslösheten	unemployment,
verktyg	tools,
barndom	childhood,
life	life,
café	coffeehouse,café,
snittet	the intersection,
huvudstäder	capital cities,capitals,
ändrade	changed,
arkiv	archive,
närvarande	present (-ly),present,
dave	dave,
kometer	comets,
övergripande	over arching,general,
chili	chili,
parterna	parties,
intag	intake,
slutliga	evenutal,ultimate,
frankrikes	frances,
castro	castro,
klarade	made it,
organisera	organize,organizing,
kontraktet	the contract,
tintin	tintin,
k	k,
brister	inabilities,
gärna	i'd love to,readily,
stämma	sue,
player	player,
tänkare	thinker,
australia	australia,
slag	kinds,
tät	compact,frequent,
serbisk	serbian,
tillhandahåller	provides,
vrida	turn,
foton	photos,
omkring	surrounding,about,around,
agnetha	agnetha,
european	european,
klimatet	climate,the climate,
josef	josef,
topp	top,
värde	value,
emi	emi,
tunn	thin,
funktioner	functions,
synder	sins,
tung	heavy,
obligatoriskt	obligatory,
finska	finnish,
lucas	lucas,
kampanj	campaign,
centraleuropa	central europe,
gudinnan	goddess,the godess,
misslyckade	failed,
manteln	the mantle,mantle,
snö	snow,
köra	drive,
koloniseringen	the colonization,
capitol	capitol,
dödsoffer	casualty,death victim,
biskop	bishop,
körs	driven,running,being driven,
birmingham	birmingham,
utrotning	extinction,extermination,
kommunal	municipal,
döda	dead,
matteus	matthew,matteus,
han	he,
vetenskapsmän	scientist,scientists,
bnp	gdp,gnp,
fysikaliska	physical,
muhammeds	mohammed's,muhammed's,
huvud	head,
hette	named,
lunginflammation	pneumonia,
har	has,have,
hat	hatred,
hav	ocean,
präst	priest,
inne	in,
underliggande	underlying,
svensson	svensson,
narkotika	narcotics,
livsstil	life style,lifestyle,
dagar	says,days,
uppmärksammade	observed,noted,noticed,
county	county,
bobby	bobby,
sedlar	bills,
alice	alice,
kust	coast,
residensstad	city of residence,county seat,
sebastian	sebastian,
ola	ola,
företräder	representing,
people	people,
parlamentarisk	parliamentary,
delade	shared,divided,split,
kulmen	the acme,peak,
fot	foot,
varierande	varying,
angränsande	adjoining,adjacent,
utser	chooses,appoints,
utses	appointed,
akademi	academy,
idéer	ideas,
myndigheter	authorities,
annan	another,
neptunus	neptunes,neptune,
stefan	stefan,
påminner	reminds,
hörde	heard,
binder	tie,
olympiska	olympic,
möjligheterna	possibilities,the possibilities,
myndigheten	the authority,
annat	other,other; another,
evangelierna	the gospels,
army	army,
o	oh,
mynnar	opening,
klubben	club,
stjärna	star,
misstänkt	accused,suspect,suspected of,
nixon	nixon,
tillverkare	producer,manufacturer,
hänt	happened,
delvis	partly,partially,
psykiska	psychic,mental,
marshall	marshall,
som	as,which,
sol	sun,
lagliga	legal,
son	son,
psykiskt	psychic,
delarna	the parts,
artikeln	the article,
hantera	handle,
nova	nova,
säkerhetspolitik	safety policy,security policy,
homo	homo,
 miljoner	millions,millon,
jönköpings	jönköpings,
offer	victim,
öppen	open,
förhållandet	relationship,
förhållanden	n/a,
öppet	open,
verde	verde,
tigern	tiger,the tiger,
avsevärt	substantially,considerably,
förväntningar	expectations,
drabbat	affected,
gymnasiet	high school,gymnasium,
drabbar	affect,troubles,afflict,
polska	polish,
syften	purpose,
pest	plague,
syftet	purpose,
fansen	the fan,
moderna	modern,
föregångare	predecessor,
konung	king,
lunds	lund's,
låtar	songs,
modernt	modern,
krävde	demanded,
ericsson	ericsson,
astronomiska	astronomical,
huvudperson	main person; main character,main character,
dotter	daughter,
aristokratin	the aristocraty,
protester	protests,
läste	read,
republik	republic,
roll	role,
olja	oil,
reggae	reggae,
avskaffades	was abolished,abolished,
bostadsområden	housing,residential areas,
jamaicanska	jamaican,
blått	blue,
vintrarna	the winters,winters,
modell	model,
transporter	transports,
danske	danish,dane,
aragorn	aragorn,
tävling	competition,contest,
noga	carefully,
sällan	seldom,rare,
povel	povel,
laddade	charged,
perioden	period,time,
kategorifödda	category: born,
förtjust	delighted,
trettio	thirty,
perioder	periods; episodes,
time	time,
erkända	acknowledged,
skatt	tax,
erkände	confession,acknowledged,
oss	us,
ost	cheese,
uppgifter	information,tasks,
stödjer	supports,
avalanche	avalanche,
uppgiften	the task,
atombomben	atom bomb,the nuclear bomb,
stålgemenskapen	steel community,
inkomst	income,
behåller	keeps,
machu	machu,
fängelset	prison,
intresserade	interested,
grön	green,
vem	who,
framställa	represent; depict; produce,produce,
marocko	morocco,marocco,
bosnien	bosnia,
musikstilar	music genres,
individer	individuals,
choice	choice,
individen	the individual,individual,
framställs	is depicted,
skillnaderna	the differences,
linné	linneus,
initiativ	initiative,
lägre	lower,
inhemska	native,
saab	saab,
oppositionen	opposition,
team	team,
uppskattningsvis	approximately,an estimated,
årig	year old,
jämnt	even,evenly,
scen	scene,
jämna	even,
firandet	celebrate,the celebration,
måne	moon,
greve	earl,
elton	elton,
köp	purchase,
kunskapen	the knowledge,knowledge,
beskydd	protection,
axel	axel,
bosatte	settled,
kön	gender,
kunskaper	knowledge,
bosatta	settled,
kusten	the coast,
katter	cats,
gula	yellow,
provinserna	provinces,the provinces,
galileo	galileo,
skydd	protection,
budskapet	the  message,the message,message,
katten	the cat,cat,
huvudsakliga	main,
studien	the study,
genomgående	consistently,pervading,
hälft	half,
landslag	national team,
studiet	the study,
studier	studies,
engelske	british,the english,english,
styrkan	strength; unit; force,strength,
publicera	publish,
kommit	to be,come,
presenterade	presented,
sprids	spreading,spreads,
samlat	single,gathered,
samlar	collect,salmar,
positiva	positive,
änglar	angels,
vuxna	adult,
sprida	spread,
judarna	jews,
positivt	positive,
samlag	intercourse,
effektiv	effective,
ställt	put,set,
dagars	day's,days,
hår	hair,
tillträdde	assumed,
ställe	place,
hål	hole,
ställa	make,set,
tabellen	the chart,table; list,
grönt	green,
straffet	the punishment,
kunskap	knowledge,
gröna	green,
påvisa	prove,
stigande	rising,
locka	attract,tempt,
missförstånd	misunderstanding,
locke	locke,
släktskap	relationship,kinship,
inkluderade	included,
rädda	save,
kretsar	circuits,circles,
utnyttjade	used,
drama	drama,
milda	mild,
årligen	yearly,
skikt	layers,
svenskan	swedish,the swede,
trigonometriska	trigonometric,
européer	europeans,
riksdagen	the parliament,
gigantiska	gigantic,
kungens	the king's,
löpande	running,assembly,conveyor (belt),
svart	black,
nyligen	recently,
data	data,
epost	e-mail,email,
portugisiska	portuguese,portugese,
stress	stress,
natural	natural,
bergarter	rock types,minerals,rocks,
undervisning	education,
påstod	claimed,
ss	ss,
sr	sr,
sv	south west,
vikt	weight,
st	saint,
sk	so called,
sm	s-m,swedish championship,
sa	said,
vika	fold,
se	see,
resulterar	result,results,
allvarliga	serious,
resulterat	resulted in,
professorn	the professor,
kong	(hong) kong,kong,
antingen	presumably,
allvarligt	serious,
clinton	clinton,
irländsk	irish,
torg	square,
ingvar	ingvar,
dialekter	dialects,
utsätts	exposed,
jim	jim,
tilldelats	awarded,
begrepp	concept,
museu	museum,
faderns	the father's,
monopol	monopoly,
personlig	personal,
hos	in; with,with,
änden	end,
öppnades	were opened,was opened,opened,
äldste	eldest,
musiken	the music,
äldsta	oldest,
matcher	games,
nation	nation,
matchen	the game,
kategoripersoner	category of persons,
kantoner	cantons,
kravet	the demand,
twilight	twilight,
musiker	musicians,
atmosfär	atmosphere,
lockar	attracts,
förväxlas	mixed up (with),confused,mistaken,
sidor	pages,
säga	say,
skivkontrakt	record contract,
dominerar	dominates,
domineras	dominated,
runstenar	runestones,rune stones,
sägs	said (to be),said,
dominerat	dominated,
födelsedag	birthday,
prisma	prism,prisma,
dynamiska	dynamic,
greker	greek,greeks,
delstaterna	states,
förstöra	destroy,ruin; destroy,
väljas	elected,be elected,choose,
hinduer	hindu,
krav	requirement,demands,
kött	meat,
riktigt	real,right,
bly	led,lead,
specifikt	specifically,
sjuka	sick,
densitet	density,
riktiga	real,
bränder	fires,
internet	internet,
roterar	rotates,
bla	among others,
sfären	sphere,
garantera	guarantee,
vård	nursing,
våra	our,
singlar	singles,
sålde	sold,
bytt	traded,switched,
byts	replaced,
väster	west,
vårt	our,
kolonier	colonies,
dramaten	dramaten,
byte	change of,
byta	switch,change,trade,
föreställning	performance,
pund	pound,
artister	artists,
punk	punk rock,punk,
flandern	flanders,
massiva	massive,
artisten	the artist,
gordon	gordon,
främst	foremost; primarily; chiefly,primarily,
givits	given,
förmån	advantage; in favor of; benefit,
hård	diffcult,hard,
potter	potter,
tsunamier	tsunamis,
hårt	hard,difficult,
open	open,
ont	bad,
urin	urine,
city	city,
tekniska	technical,
flytande	floating,liquid,
teologi	theology,
skådespelarna	actors,
råolja	crude oil,
intill	beside,adjacent to,
sjö	naval,lake,
nästa	next,
williams	williams,
animerade	animated,
vilka	who; which; that,who,
tillräckligt	sufficient,
irakiska	iraqi,irakish,
tillräckliga	sufficient,
svenskarna	the swedes,
yttersta	furthest,supreme,highly,
provins	province,
dygn	day,
fiskar	fishes,
uppenbarelser	revelations,
berlinmuren	berlin wall,the berlin wall,
kamprad	kamprad,
motståndarna	the opponents,opponents,
tankar	tank,thoughts,
sak	thing,matter; case,
san	san,
generation	generation,
konsekvenser	consequences,
argument	argument,
församlingar	parishs,
känslan	feeling,the feeling,
burundi	burundi,
allen	allen,
utgåva	edition,issue,
staden	city,the city,
priserna	prices,the prices,
övriga	other,
takt	rate,
ambassad	embassy,
zon	zone,
jefferson	jefferson,
massa	mass,
övrigt	other,
förändringen	the change,
föder	give birth,gives birth,give birth of,
muslimer	muslims,
finlands	finland's,finlands,
sekreterare	secretary,
knep	tricks,sleight of hand,
religionen	religion,the religion,
betyda	mean,
religioner	religions,
forskningen	the science,
driva	operate,run,
frihetliga	libertarian,
inledningen	introduction,
ursprung	origin,root,
rykte	reputation,
sades	said,was said,
drivs	driven,
rött	red,
olagligt	illegal,
axl	axl,
genomförts	out,
beckham	beckham,
dimensioner	dimensions,
ormar	snakes,
sjöss	sea,
antalet	number,the number,
stärkte	strengthened,increased,
slog	hit,
hockey	ice hockey,hockey,
beatles	beatles,
katoliker	catholics,
platta	flat,
undersöka	research,
rörande	concerning,
spetshundar	tip of dogs,
ländernas	the countries,countries',
artist	artist,
råd	advice,council,
översättningen	translation,the translation,
roger	roger,
ledningen	the lead,
ljudet	the sound,
varna	varna,
yta	surface,
monark	monarch,
erbjöds	offered,
dagsläget	present situation,
hämtar	is,gets,
spetsen	edge; top,tip,
brännvin	schnaps,
snabbare	faster,
behovet	need,the need,
nederbörden	the precipitation,
skärgård	archipelago,archipelagos,
talman	spokesperson,president,speaker,
personlighet	personality,
enhetlig	unitary,uniform,
utgörs	consists of,make up,
förvaltning	administration,
källa	source,
kritiserade	critisized,criticized,criticised,
begränsningar	limitations,
upplever	experience,
kontrakt	agreement,contract,
utgöra	compose,make up,
kilometer	kilometer,kilometers,
revolutionär	revolutionary,
små	small,little, small,
gäller	of,refer to,
amerikanskt	american,
anledningarna	reasons,the reasons,
söka	search,
screen	screen,
fynd	finding; finds,
antika	ancient,
amerikanske	american,the american,
jobb	job,
amerikanska	american,
galaxer	galaxies,
basisten	basist,the basist,
skönlitteratur	fiction,
mans	man's,
erics	erics,
rekord	record,
mani	mani,mania,
tillsätts	appointed,appoints,
upproret	the upprising,revolt,
klimat	climate,
hamnade	landed,ended up,
anta	assume,assume; adopt,
drogs	was pulled,
farfar	paternal grandfather,
bolag	company,
luft	air,
cupen	the cup,
lidit	suffered,
formen	the form,
formel	formula,
sångerska	songstress,singer,
warhol	warhol,
tillåter	allows,allow,
tillåtet	allowed,
pernilla	pernilla,
former	forms,
landskapen	the landscapes,landscape,
samling	collection,
vojvodina	voyvodina,
landskapet	landscape,
friska	healty,
situation	situation,
föregångaren	predecessor,it's predecessor,
peruanska	peruvian,
aborter	abortions,
aluminium	aluminum,
startar	begins,
bror	brother,
ekonomi	economy,
tillåtelse	permission,allowed,
sammanfaller	coincides,
ohälsa	disorders,
världsbanken	world bank,
undersökning	survey,
träffat	met,
ärftliga	genetic,
otto	otto,
träffas	meet,
oceanen	the ocean,
ekologi	ecology,
nationalparker	national parks,
singapore	singapore,
sägas	is said,is said (to be),
lindgrens	lindgren's,lindgrens,
förkortning	abbreviation,
senator	senator,
dsmiv	dsm-iv,
personlighetsstörning	personality disorder,
costa	costa,
tillfälle	instance,occasion,
gestalter	beings,figures,
avser	regards,regard,
avses	refered,regard,referred,
ifrågasatt	questioned,
iraks	iraq,
summer	sommar,
förluster	losses,
bokförlaget	bokförlaget,publisher,publishing house,
berättelse	tale,
rest	remain,rest,
koncentration	concentration,
spårvagnar	trams,
psykologisk	psychological,
likheter	similarities,similarity,
resa	travel,
libyen	libya,
förlusten	loss; defeat,
judarnas	jews,
kastar	throws,to throw,
heliga	holy,holy; holy,
unika	unique,
sprider	spreads out,spread,spreads,
helige	holy,
miljon	million,
instrument	intrument,
körberg	körberg,
sänka	lower,
infördes	introduced,
unikt	unique,
heligt	holy,
snart	soon,
vinkel	angle,
dark	dark,
jorderosion	earth erosion,soil erosion,
unesco	unesco,
litteraturen	literature,
skadade	wounded,damaged,
stammar	tribes,
statsreligion	state religion,
vattenånga	steam,water vapour,
carl	carl,
ekonomier	economies,
stupade	fallen,killed,
fossila	fossilized,
intet	nothing,
jobbar	work,does the work,
nämnas	mentioned,worth mentioning,
domkyrkan	the cathedral,
ursprungsbefolkning	native population,
kännedom	knowledge,
inkluderas	is included,
björn	björn,
föreslog	suggested,propose,
institutionerna	institutions,
än	than,yet,
exil	exile,
cannabis	cannabis,
varsin	(one) each,
atomkärnor	nuclear particles,atomic cores,
västerås	västerås,
katolsk	catholic,
jacksons	jackson's,jacksons,
medlemsstater	member states,member-state,
organisationen	organization,the organization,
herrlandslag	men's national team,
vissa	some,
populationen	the population,
befinner	placed; situated; positioned; are,
digerdöden	the black death,
populationer	populations,
wien	vienna,
organisationer	organisations,
industri	industry,
visst	certain,
regissör	director,
berger	berger,
upplevelser	experiences,
berget	the mountain,
image	image,
partiet	the party,
partier	parties,
angola	angola,
bergen	the mountains,mountain,
het	up to date,
striderna	the battles,
förintelsen	the genocide,
philadelphia	philadelphia,
evangeliska	evangelical,
söker	searches,seek,seeks out,
hel	(whole) lot (of),
hamnen	the harbour,
sover	sleep,
mediet	the medium,
hänger	depends,
hänvisning	reference,
hells	hells,
bevarat	preserve,preserved,
bevaras	are protected,
mick	mick,mike (microphone),
utvecklandet	development,
existerande	existing,
bevarad	kept,preserved,
åttonde	the eighth,
rush	rush,
sällskap	company,
jamaicas	jamaicas,jamaica's,
hexadecimalt	hexa-decimal,
kvartsfinalen	quarter finals,quarterfinals,
utmed	along,
vinkeln	the angle,
afrodite	afrodite,
förbundsstat	federal,federal state,
produkt	product,
puls	pulse,
krona	crown,
ac	ac,
brodern	the brother,
johnny	johny,
redovisas	shown,accounted for,
gustafs	gustafs,gustaf's,
am	am,
al	alder,
bronsåldern	bronze age,the bronze age,
beordrade	ordered,
övernaturliga	supernatural,
håll	ways,
väsentligt	substantially,relevant,
testamentet	testament,
vore	would,
truman	truman,
federala	federal,
rökning	smoking,
innehåll	content,
belönades	rewarded,awarded,
svåra	difficult,
avslöjade	revealed,
såsom	like,
gifta	marry,
värmlands	värmlands,
koppar	copper,
gifte	married,
medverkan	the contribution,
kvarstod	remained,
medverkat	participated,
värd	worth,
terry	terry,
vanliga	ordinary,regular,usual,
forntida	prehistoric,
kommunen	municipality,
kommuner	counties,
beteckning	indication,label,
adam	adam,
omgivningen	surroundings,the surrounding,
decennierna	decades,the decades,
original	original,
renässans	renaissance,
känslor	feelings,
släppt	released,relinquished,
släpps	(is) released,
elektron	electron,
halsen	the neck,the throat,
anpassning	adaption,
kammare	chamber,
års	years (age),years,
släppa	release,
likartade	similiar,similar,
 kmh	km/h,
norr	north,
skogarna	the forests,forests,
pojkvän	n/a,boyfriend,
ullevi	ullevi,
tv	tv,
romanen	novel,
nederbörd	precipitation,
mildare	cooler,milder,
romaner	novels,
th	th,
nord	north,
te	tea,
angående	concerning,
ta	take,
avlägsna	distant,remove,
använder	using,uses,
arvet	the inheritance,
telefonen	the telephone,
strand	beach,
utländsk	foregin,foreign,
sant	true,
ensamma	alone,
djurarter	species of animals,animal species,species,
borrelia	borrelia,
muslimska	muslim,
utsåg	declared,
sand	sand,
siffrorna	the numbers,numbers,
områdets	the area's,of the area,
harry	harry,
sann	true,
språkbruk	language (use); parlance; phraseology,parlance,
förmedla	pass; express; mediate,
döttrar	daughters,
samoa	samoa,
påståenden	claims,assertions,
synd	sin,
dödsstraff	death penalty,
utökade	expanded,increased,
pass	an,
givaren	donor,the giver,dealer,
syns	seen,
richard	richard,
delen	part,
soldater	soldiers,
islams	islams,islam's,
leif	leif,
gjorts	done,
hänsyn	consideration,
full	full,
gruppen	the group,
själen	soul,the soul,
arkeologiska	archaeological,
november	november,
legend	legend,
motstånd	resistance,
äventyr	adventure,adventures,
hindra	prevent,
traditionella	traditional,
exklusiv	exclusive,
traditionellt	traditional,
social	social,
action	action,
oftare	more often,
varelser	creatures,
sena	late,
kommunistpartiet	the communist party,
vid	in,by,at,
ordinarie	permanent,ordinary,regular,
vii	vii,
vin	whine,wine,
juridiskt	juridical,
vis	wise,
kuiperbältet	the kuiper belt,the cuyper belt,
vit	white,
främja	further,promote,
skapa	create,
biskopen	the bishop,
mors	mothers,
petroleum	petroleum,
underordnade	subordinates,
pearl	pearl,
sitter	serve,
presenterades	presented,
rhen	the rhine,
dödligt	lethal,deadly,
mora	mora,
fyrtio	forty,
bevis	evidence,
mord	murder,
ragnar	ragnar,
uppskattad	estimated,appreciated,
berättade	told,
uppskattas	is appreciated,appreciated,
graven	the grave,
schweiz	switzerland,
undergång	during navigation,doom,destruction,
socialt	social,
inträffade	occurred,happened,
medelklassen	middle class,
science	science,
beskyddare	protector,
monoteistiska	monotheistic,
cykel	bicycle,
morgan	morgan,
kapitalism	capitalism,
studenter	students,
läkaren	the doctor,
samväldet	the commonwealth,
jakob	jakob,
säljas	is sold,
nordvästra	northwest,north western,
skadliga	harmful,
staten	state,
mellersta	middle,the middle,
drabbades	affected,where hit by,afflicted,
spansk	spanish,
järnvägsnätet	railroad network,
information	information,
vägnätet	road network,
hugo	hugo,
uppfattade	perceived,perceive,
ansetts	regarded,regarded; viewed (as),
uppnått	met,achieved,
lejon	lion,
riksdagens	the parliament's,the parliaments,
retorik	rhetoric,
brett	broad,
kedjan	the chain,
produktionen	the production,
referens	reference,
lanka	lanka,(sri) lanka,
köpte	bought,
barnens	the child's,childrens,
komplext	complex,
anklagade	accused,
pucken	the puck,
komplexa	complex,
utvidgning	enlargement; expansion,
hållit	held,maintained,kept,
nationerna	the nations,nations,
aktiviteten	the level of activity,
östblocket	east block,the eastern bloc,
scott	scott,
kvinnors	women's,
aktiviteter	activities,
anställda	employed,
radion	the radio,
känsla	feeling,
alla	all,everyone,
högskola	college,
protestanter	protestants,
caesars	caesars,
termen	the term,term,
termer	term,
alls	all,
få	have; make; few,
stadshus	town hall,city hall; town hall,
isaac	issac,
konstruerade	constructed,
samhällets	of society,
känner	know,
källan	source,the source,
beräkna	calculated,calculate,
privilegier	privileges,
inledande	initial,
produceras	produced,
producerar	produces,
grekisk	greek,
producerat	produced,
introducerade	introduced,
producerade	produced,
olycka	accident,
intåg	entry,advent,
budskap	message,
målning	painting,
blodet	the blood,
denne	that he,
genom	through,
härrör	derived,
enstaka	occasional,single,
england	england,
populärt	popular,
sydöst	south east,
populära	popular,
blues	blues,
förespråkade	advocate,
kretsen	the order,
finner	finds,
uppfördes	was constructed,constructed,
massiv	massive,
omröstningen	the election,
kopplad	connected to,connected,
garvey	garvey,
avgick	resigned,retired,
norska	norwegian,
uppstått	arised,arisen,
sammanfattning	summary,
besökte	visited,
kopplat	coupled; connected,connected,
hallucinationer	hallucinations,
medel	middle,
sparken	gets fired,fired,
alltmer	increasingly,more and more,
stjärnor	stars,
driver	drive,
båda	both,
både	both,
kostade	cost,
ålands	Åland island's,the Åland island's,
kärnkraft	nuclear power,
poeten	the poet,
teknologi	technology,
definition	defined,definition,
service	service,
turistmål	tourist destination,tourist attraction,
gatorna	the streets,
naturens	nature's,
omfattar	encompass,
skolan	school,
w	w,
nivåer	levels,
besök	visit,
uppenbarelse	apparition,revelation,
principen	the principal,
bidragit	contributed,
kristna	christian,
foten	foot,
skiftande	shifting,
spekulationer	speculation,speculations,
såg	saw,
gemensamma	common,
avel	breeding,breed,
liknas	compared to,likened,
liknar	similar to those,
saint	saint,
sår	wound,
besläktat	related to,related,
läggas	laid,added,
chefen	commendant; commander,
tappade	lost,
zeus	zeus,
zeppelin	zeppelin,
moder	parent,mother,
svår	difficult,
grace	grace,
obama	obama,
organiseras	organizes,
återkom	returned,
niklas	niklas,
marknadsekonomi	market economy,
organiserad	organized,
nikolaj	nikolaj,
ägg	egg,
äga	own,
väljer	elects,
avslutade	ended,
inkluderar	includes,
generationen	generation,the generation,
inkluderat	included,including,
ägt	taken,
generationer	generations,
astronomin	the astronomy,
visats	shown,
framåt	forward,forth,
varianten	version,variant,
norstedts	norstedt's,norstedts,
without	without,
varianter	variants,diversities,
vinterspelen	winter games,
arabisk	arabic,
edison	edison,
sydostasien	south east asia,
brooklyn	brooklyn,
plan	level,
kombinationer	combinations,
arter	species,
utsattes	subjected,were exposed,
cover	cover,
kanalen	the channel,
kanaler	channels,
förklaringen	the explanation,
kombinationen	the combination,combination,
golf	golf,
omfattade	covered,
pengarna	the money,
presidentens	the president's,the presidents,
detalj	detail,
karaktär	character,
falskt	false,
richmond	richmond,
framgångar	success,
existensen	existence,
betydelser	meanings,
jämföra	compare,
befolkningstätheten	n/a,
wayne	wayne,
betydelsen	the meaning,
jämfört	compared,compared (to),
kontor	office,
karakteristiska	characteristic,
genomgick	underwent,
gratis	free,
evolutionen	the evolution,
tekniken	techinque,the technology,
tekniker	technician,
utbildningen	education,
föll	fell,
erkännande	recognition,
victoriasjön	lake victoria,
tanken	the thought,idea,
ledare	leader,
bytet	the exchange,
populärmusik	popular music,pop music,
byten	byte,
kill	kill,
anslutning	connection,
sköt	shot,
någon	someone,
kriterier	criteria,
ses	are seen,
ser	see,sees,
koranen	the koran,the quran,
sex	six,
sed	thirst,
psykologiska	psychological,
uppkomsten	origin,
märta	märta,
järnväg	railroad,railway,
sen	since,
något	something,
sorters	kinds,
institutet	institute,the institution,
församlingen	parish,congregation,
påverkat	influenced,
guinea	guinea,
neutralitet	neutrality,
fission	fission,
stärkelse	starch,
alqaida	al-qaida,al-qaeda,
rita	paint,draw,
europe	europe,
europa	europe,
giftermål	marrige,marriage,
medveten	conscious,aware,
avvikelser	deviations,derivations,
stadsdel	city district,neighborhood,district,
demografiska	demographic,demographical,
forskare	researcher,scientists,
bästa	the best,best,
medicinering	medication,
förändring	change,
bäste	best,
messias	messiah,
stå	stand,
halmstads	halmstad's,
kopia	copy,
samma	the same,same,
transeuropeiska	trans-european,transeuropean,
upprättades	establish,
krisen	the crisis,
kriser	crises,
luis	luis,
allierade	allied,allies,
decennium	decade,
sommaren	summer,the summer,
koalition	coalition,
mått	measure,
väntade	expected,expected; were waiting,waited,
tillväxt	growth,
potentiellt	potential,
kyrilliska	cyrillic,
idén	the idea,
blod	blood,
pågår	(in) progress,
föranledde	brought about,led,
beskrevs	was described,described,
skönhet	beauty,
östafrika	east africa,
fira	celebrate,
hovrätten	the court of appeal,
fritz	fritz,
uppleva	experience,
fritt	free,
föreningar	associations,organizations,
systematik	systematics,systematic,
handling	act,
framträder	appear,stand out,
projekt	project,
budget	budget,
guldbollen	guldbollen,
individerna	the individuals,
bestående	lasting,
brottslighet	criminality,crime,
pressen	the pres,
real	real,
arbete	work; labor,
von	von,
motors	engine's,
teoretisk	theoretical,
erkänna	recognize,
lokaler	studios,place,
korruptionsindex	corruption index,
hovet	court,the court,
kritiker	critics,critiques,
barney	barney,
möjlighet	an opportunity,oppertunity,possibility,
omvandlas	convert,converted,
omvandlar	transmuted,
skalet	shell,the shell,
högste	supreme,highest,
barnen	children,
arméer	army,
kritiken	the criticism,the critique,
laddning	charge,
centrum	center,
debatter	debates,
republiken	the republic of,the republic,
republiker	republics,
debatten	debate,the debate,
kring	around,
djurgården	djurgården,
vargar	wolves,
euro	euro,
normala	normal,
phil	phil,
krigsmakt	military power,armed forces,
person	person,
kontakter	contacts,
konkret	concrete,
tunnelbana	subway,
stränder	beaches,
släppas	released,be released,
telegram	telegram,
stockholms	stockholm's,
finansiella	financial,
kontakten	the contact,
mandat	mandate,
fascistiska	fascist,fascistic,
relationer	relations,
festivalen	festival,the festival,
tobak	tobacco,
nordväst	north west,northwest,
festivaler	festivals,
jönssonligan	jönssonligan,
tomas	tomas,
hennes	her,
format	shaped,format,
kopplas	connected,
turnéer	tours,
melker	melker,
avvisar	reject,
skara	city in south-central sweden (uppland),crowd,
samarbete	collaboration,
ivar	ivar,
västsahara	western sahara,
samarbeta	cooperate,
da	da,
talrika	numerous,
funnit	found,
skarp	sharp,
utlösa	trigger,
informationen	the information,
patrick	patrick,
ivan	ivan,
alexandra	alexandra,
ulrich	ulrich,
lenin	lenin,
saknar	lacks,lack(-s),missing,
saknas	missing,
användbar	useful,
utvecklades	(was) developed,
avskaffade	abolished,absolished,
saken	the thing,the matter,
ovan	above,
wallenstein	wallenstein,
öka	increase,
brasilianska	brasilian,
trafiken	the traffic,
turnerade	toured,
religion	religion,
riksförbundet	national association,
säger	says,claims; says,
nybildade	newly formed,newly established,
tåg	trains,
ugandas	of uganda,
västra	west,
bl	short of "bland" - in the context: bl. a (bland annat) = among others,
vagnar	wagons,carriges,
bo	living,
plocka	pick,
engelska	english,
bokstav	letter,
santa	santa,
by	village,
ideologin	ideology,the ideology,
bosättningar	settlements,
soldaterna	soldiers,the soldiers,
dagligen	daily,
aggressiv	aggressive,
arméerna	armies,
stuart	stuart,
fungerande	effective,working,
papper	paper,
inte	not,
inta	taken,
colorado	colorado,
syret	the oxygen,
hemingway	hemingway,
efterföljande	subsequent,
spridas	spread,
kraven	the demands,requirements,
popsångare	popsinger,pop singer,
uppkallad	named,
producent	producer,
förlaget	publisher,the publisher,the publishing company,
seger	victory,
veckor	weeks,
utbröt	erupted,broke out,
samerna	the lapp,
knuten	tied to,bound,
hälften	the one half,half,
fattigdom	poverty,
förbindelse	connections,
begreppen	the concepts,the terms,
söder	south,
rörlighet	movement,
pastor	pastor,
begreppet	term,concept,
posten	the position,
atom	atom,
kritisk	critical,
lovade	promised,
lina	line,lina,
dröm	dream,
fader	father,
cia	cia,
ut	out; up,out,
dom	judgement,conviction,
drogmissbruk	drug abuse, substance abuse, drug addiction,
up	up,
us	oss,
ur	from,out,
konventionella	conventional,
distrikt	district,
uk	uk,
protestantiska	protestant,protestantic,
inriktade	oriented,
testamente	will,wills,
professor	professor,
översvämningar	floodings,
nämner	mentions,
dog	died,
diverse	some,
utbyggt	develpoed,built,extended,
makedonska	macedonian,makedonish,
nationalism	nationalism,
inblandning	involvement,incorporation,
matematiken	mathematics,
händelsehorisonten	event horizon,the event horizon,
räkna	count,
värld	world,
edwards	edward's,
skrivits	been written,
innehåller	include,contains,
nordafrika	north africa,
innehållet	content,contents,
matematiker	mathematician,
siffror	numbers,
upplaga	edition,submission,
individuella	individual,
besegra	defeat,
dominerades	was dominated,
radikala	radical,
djurgårdens	djurgården's,
ägnar	spend time,dedicated,
grovt	heavy,roughly,
riskerar	risks,there is a risk,
springsteen	springsteen,
radikalt	radical,radically,
slås	beat,is hit,
alltså	so,therefore,really,
land	country,
passagerarna	passengers,the passengers,
uppträdande	performance,appearance,
symtom	symptom,
age	do,age,
härstammar	derived,stems,
sawyer	sawyer,
texter	texts,
inspelning	recording,
persbrandt	persbrandt,
släpptes	was released,
alltför	all too,exessive,
bakåt	reverse,
anorektiker	anorectics,
turkisk	turkish,
dyraste	most expensive,
hamnar	lands,ports,
hamnat	got,ended up,got in to,
listade	listed,
dickinson	dickinson,
dancehall	dance hall,
sent	late,
lärde	learned,
märken	brands,sign,
hustru	wife,
palestinier	palestinians,palestinian,
kommunistiska	communistic,communist,
drogen	the drug,
berömda	famous,
överleva	survive,
tillhörande	belonging to,belonging (to),
magic	magic,
tro	think,
påverka	influence,
eva	eva,
tre	three,
jobbet	the job,
romerska	roman,
överlevt	survived,
romerske	roman,
opinionen	opinion,
leonardo	leonardo,
bolsjevikerna	the bolsheviks,
regelbundna	regular,
ställde	stood up,
årtionden	decades,
förhållandevis	relatively,
förkortningar	abbreviations,
pris	price,prize,
antog	adopted,
index	index,
expressen	expressen,
indiens	india's,indias,
suveräna	terrific,supreme,sovereign,
möjliggör	enables,
birk	birk,
indian	indian,
ledande	leading,
wembley	wembley,
stadskärna	city core, city center,town centre,
led	suffered,
lee	lee,
lyckades	succeeded,
sålunda	thus,
leo	leo,
lev	live,
hälsa	tell (him i said hi),
talang	talent,
begravd	buried,
motorvägarna	the highways,
casino	casino,
titanic	titanic,
anländer	arrive,arrives,
tillkom	resided,
insulin	insulin,
högsta	highest,
opinion	opinion,
huvudvärk	headache,
emot	against,
förlora	lose,
oxenstierna	the oxenstierna,
mening	sentence,
indianerna	the indians,
anatolien	anatolia,
andreas	andreas,
varmare	warmer,
rico	rico,
elever	students,
godkänna	approve,
klaviatur	keyboard,
toy	toy,
orkester	orchestra,
existerade	existing,
författning	constitution,
samspel	interaction,teamwork,
ytterst	very; extremely,highly,
överlevande	survivor; survivors; surviving,
villor	houses,villas,
edwall	edwall,
lokalt	locally,local,
nordliga	northernly,northern,
advokat	lawyer,
lokala	local,
peka	point (at; to; in),point,
sekel	century,
upprätthålla	maintain,keep up,
process	process,
klassisk	classic,
etta	number one,
syre	oxygen,
high	high,
tryckta	printed,
sydöstra	the southeast,south east,south eastern,
föregående	preceeding; previous,previous,
halmstad	halmstad's,
gitarr	guitar,guitarr,
saknade	lacked,missed,
delad	divided,
övergrepp	assault,abuse,assult (-s),
hormoner	hormons,
delas	shared,
delar	proportions,parts,
delat	divided,
sydvästra	southwest,
kriminella	criminal,
gunwer	gunwer,
amerika	america,
djurens	the animals,
profeten	the prophet,
profeter	prophets,profets,
regeringsmakten	govermental power,government power,
platt	flat,
väckt	awaken,woken,
slutsatser	conclusions,
frågor	questions,
lundgren	lundgren,
nancy	nancy,
napoleons	napoleon's,
byggnadsverk	building,
borde	should,
handboll	handball,
diskar	disks,
möjligt	possible,
hårdast	the most,
universiteten	universities,the universities,
frånvaro	absence,
hunnit	reached,had,had time to,
universitetet	the university,
bensin	gasoline,
möjliga	possible,
solvinden	the solar wind,solar wind,
västerbottens	västerbotten's,
eliten	the elite,
uppdelat	divided,split,
fristående	independent,stand-alone,
tecknet	the sign,sign,
uppdelad	split,
puerto	puerto,
beståndsdelar	elements,
ovanlig	unusual,
bekant	known,acquaintance,
bryter	breaks,breaking; violating,
hemmaplan	home,home turf; domestic (level),
dock	however,
kiss	kiss,
rotation	rotation,
huvuddelen	main part,
sönder	broken,
symboliserar	symbolized,
peking	beijing,
välfärd	wealth,
intressen	interests,
fortsätta	continue,
smallwood	smallwood,
överföras	transferred,
astronomer	astronomers,astronomer,
intresset	interests,the interest,
bay	bay,
etymologi	etymology,
matrix	matrix,
olika	different,
trycktes	was published,
utbildad	educated,
enskilda	individual,
anledningen	reason,
umgänge	company,
kapitalismens	capitalism's,
marxistiska	marxist,
bekräftades	confirmed,was confirmed,
fram	until,
undertecknades	signed,
redskap	device,
högtid	festival,festival; holiday,
mötte	motte,met,
kalle	kalle,
påverkats	influenced,affected,
underverk	wonder,
uppe	up,(on) top, up, above,
lundin	lundin,
förts	brought,
tempererat	temperate,tempered,
dubbel	double,
liggande	placed,lie,
kompositör	composer,
krävt	taken,
våldsam	violent,
krävs	needs,required,
david	david,
blanda	mix,
krets	sphere,circuit,
helst	rather,anyone,any time,
davis	davis,
hussein	hussein,
kräva	demand,
skillnad	difference,
playstation	playstation,
åring	years,
komplicerade	complex,
jesus	jesus,
användningsområden	possible use,applications,
schweiziska	swiss,
muhammad	muhammad,
nordkoreanska	north korean,
studerade	studied,
värdefulla	valueable,valuable,
festival	festival,
system	system,
bygget	the construction,
syster	sister,
hebreiska	hebrew,
tränga	push (aside),cut in,
teatern	the theater,
blivit	become,
utbyggnad	development,addition,expansion,
pristagare	prizewinner,
konservativ	conservative,
haven	the seas,
visdom	wisdom,
hampa	hemp,
samverkar	co-operating,co-operates,
roberto	roberto,
väsen	entity,
roberts	roberts,
reagans	reagan's,
troende	faithful,
samverkan	co,cooperation,
jonatan	jonatan,jonathan,
räcker	enough,
användaren	the user,
inre	inner,
förslag	proposal,
flygplats	airport,
kritiskt	critical,
instruktioner	instructions,
lindh	lindh,
sinatra	sinatra,
sekvens	sequence,
kritiska	critical,
best	best,
linda	linda,
viss	certain,
slutsatsen	the conclusion,
när	when,
nät	web,net(work),
trosbekännelsen	faith of confession,
slovakien	slovakia,
vardagen	the weekday,
kvinnliga	female,
uppror	uprising,rebellion,
flyga	fly,
förutsättningarna	prerequisites,
medan	while,
framgår	is shown,
synliga	visible,
våren	the spring,
bred	broad,
bokstaven	the letter,
nordöst	northeast,
synligt	wisible,seen,visible,
befolkningens	population's,
brev	letter,
beteende	behaviour,behavior,
uppdelade	divided,
tyvärr	unfortunately,
hopp	hopes,hope,
fursten	prince,
östfronten	the east front,
samisk	samian,
jan	jan,
religionens	religion's,
liksom	and,as is,
jah	jah,
jag	i,
skarsgård	skarsgård,
ilska	anger,
handla	act; buy; consume,act,
abba	abba,
parlamentet	the parlament,
lägger	put,lies,add,
fotbollsspelare	football player,
generalen	the general,
bonde	bonde,farmer,
parlamenten	the parliament,
halvklotet	hemisphere,
britterna	british,the brits,
h	h,
rowling	rowling,
effekterna	the effects,effects,
iranska	iranian,
rymmer	has,holds,
guvernör	governor,
myndigheterna	authorities,the authorities,the authoroties,
debuterade	debuted,
michail	michail,
konungarike	kingdom,
avlidit	perished,died,
priset	the prize,
kronisk	chronic,
uppträdde	appeared,perform,
lämplig	suitable,
freddy	freddy,
vietnams	vietnam's,
författarskap	the writer,authorship,
sjöng	sang,
upprättandet	establishment,
längst	farthest,
sjönk	sunk,sank,
balansen	balance,the balance,
kategorisvenskar	category swedes,
striden	fight,
finalen	final,
bolivias	bolivia's,
strider	strides,conflict,battles,
bilar	cars,
ende	only,
förklaringar	explanations,
kedjor	chains,
islamiska	islamic,
ett	a,one; a; an,
marknaden	the market,
figuren	the character,figure,
religiöst	religious,
tycker	think,thinks,
fåglar	birds,
egypten	egypt,
norge	norway,
marknader	markets,
ogillade	disliked,
belägen	located,situated,
tätbefolkade	densely populated,
ekvatorn	equator,the equator,
religiösa	religious,
botten	the base,bottom,
dör	dies,
malcolm	malcolm,
mengele	mengele,
cd	cd,
sannolikhet	probability,
död	dead,
bröllop	wedding,
stabila	stable,
musikvideo	music video,
öst	east,
dök	dove,turned,
antal	number of,
jussi	jussi,
keltiska	celtic,
företaget	the company,
överallt	everywhere,overall; everywhere,
centralort	central city,regional centre,
växt	plant,
genetik	genetics,
moraliska	moral,
företagen	the companies,
antas	is required,expected (to),
antar	adopt,suppose,
typisk	typical,
frågorna	questions,questions; issues,
molekyler	molecules,
föreställer	picture,depicts,
atlanta	atlanta,
mandatperiod	term,term (of office),term of office,
långsamma	slow,
erhöll	recieved,acquire,
rikets	the realms,its,the kingdom's,
demokrati	democracy,
aktivitet	activity,
vd	ceo,
ondskan	the evil,
förlopp	pattern,developments,
omnämns	is mentioned,
vi	we,
ryssland	russia,
vm	world championship,
lust	desire,
flickor	girls,
skapare	creator,
föreligger	is,exist,
sitt	its,
referenser	references,
evenemang	event,
spela	play,
tupac	tupac,
armé	army,
känt	known,famous,side,
juan	juan,
medeltida	middleaged,medival,
huden	skin,
paulo	paulo,
matthew	matthew,
josé	jose,
känd	known,famous,
terrorism	terrorism,
flesta	most,
columbia	columbia,colombia,
sade	said,
konstantin	constantine,
framförde	presented,
anordnas	organised,arranged,
anfield	anfield,
ikea	ikea,
sjukhus	hospital,
diabetes	diabetes,
representera	represents,represent,
obamas	obama's,
mänskligt	human,
klubbarna	the clubs,
väger	weighs,weight,
vägen	the road,
mänskliga	human,
ledda	led,run (by),
uno	uno,
versaillesfreden	treaty of versailles,
mellanrum	space,
kontakt	contact,
summan	sum,the sum,
renässansen	the renaissance,
paul	paul,
pappa	dad,
tolkade	interpreted,
förknippas	associated to,associated,associate,
kunder	customer,customers,
planeter	planets,
frågan	the question,
englands	england's,
planeten	planet,the planet,
kosovos	kosovo's,
filmens	the film's,
framtid	future,
förknippad	associated,
motorvägen	motorway,highway,
ledarna	the leaders,
gul	yellow,
dess	then,its,
arbetarklassen	working class,the working class,
tillverkning	production,
pressas	pressed,
följeslagare	companion,
lät	had,sounded,
emma	emma,
lär	teach,learn,
aktiebolag	limited company; joint-stock company,stock company,
vallhund	herding dog,
stadsbild	cityscape,
amazonas	the amazon rainforest,amazonas,
symptomen	the symptoms,
högskolan	hogs school,university,college,
flotta	fleet,
uppskattades	appreciated,was appreciated,
tackade	thanked,said/thanked,
visade	showed,showed; displayed,
miniatyr|	miniature,
anarkismen	the anarkism,anarchism,
trotskij	trotskij,
lägsta	lowest,
stannar	stays,stay,
transport	transportation,transport,
skriftliga	written,
sällskapet	the company,
morris	morris,
kolonin	colony,
behandlades	treated,
toppar	tops,(that) peaks,
tänkandet	thinking,the way of thinking,
dags	time,
naturlig	natural,
kollektivtrafik	public transport,
ateist	atheist,
svaga	faint,weak,
fråga	ask,question,
biologi	biology,
ateism	atheism,
östberlin	east berlin,
svagt	weak,
smärta	pain,
vargen	the wolf,
användande	use,use; usage,
kontinenten	the continent,
må	may,
basis	basis,
höger	right,
blodiga	bloody,
angeles	angeles,
kontinenter	continents,
absint	absinthe,
hittills	so far,
burma	burma,
anpassade	custom,
släpper	releases,
upplösningen	disbandment,
sekelskiftet	the turn of the century,
planetens	the planets,
kristus	christ,
lund	lund,
mera	more,
varma	warm,
bedöma	judge; decide,
skola	school,
blå	blue,
fläckar	stain,stains and spots,
bedöms	judged,evaluated,
överbefälhavare	commander-in-chief,
tina	thaw,
förra	last,former,
samlingar	collections,
förre	former,
indonesien	indonesia,
apollo	apollo,
socialistiska	socialistic,
svält	starvation,starvations,
återkommer	returning,
volvo	volvo,
ruset	the fuddle,
stormakt	great power,major power,
monument	monument,
inrättades	established,
distribution	distribution,
butiker	shops,stores,
ovanför	over,above,
kingston	kingston,
heter	(is the) name (of),is named,
utnyttjar	uses,
utnyttjas	utilized,used,
skilsmässa	divorce,
separerade	separated,
särskild	specific,particular,
banan	the track,banana,
vitryssland	belarus,
månader	months,
sharia	sharia,
programmet	the application,the program,
öga	eye,
distinkta	distinct,
lutning	angle,incline,
relationen	the relation,
månaden	the month,
oavgjort	draw,
modernistiska	modernistic,
bröd	bread,
övergång	transition,
francisco	francisco,fransisco,
uttalade	commented; made a comment; spoke about,spoke,stated,
tider	times; ages,times,
förhandlingar	negotiations,
bröt	broke,
tiden	the time,time,
inspiration	inspiration,
syskon	sibling,siblings,
sänker	lowers,sinks,
jordbävning	earthquake,
utseende	appearance,
kommersiell	commercial,
nederländska	dutch,
brevet	the letter,
näsan	the nose,
representanthuset	house of representatives,
invadera	invade,
preussen	prussia,
konsekvenserna	consequensis,
energikälla	energy source,energy call,
barmel	barmel,
bibel	bible,bilble,
spel	game,
edward	edward,
grundande	founding,
ren	deer,
samhället	the society,society,
mördade	murdered,
stödde	supported,
golvet	the floor,
främsta	primary; foremost; primarily; principally,
främste	premier,
jacob	jacob,
skolor	schools,
special	special,
innefattar	includes,
uttryck	expression,
estland	estland,estonia,
jamaica	jamaica,
starkast	strongest,
ständerna	the cities,
sabbath	sabbath,
horn	horns,horn,
alltsedan	even since,since,
förbättringar	improvements,
eurovision	eurovision,
italiens	italy's,italian,
verksamma	active,
kraftfull	forceful,powerful,
tolv	twelve,
bidrag	contribution,
vampyr	vampire,
cyklar	bicycles,bikes,
bidrar	contributes,
petra	petra,
musikalen	the musical,
räddar	saves,saved,
bortgång	passing,
pluto	pluto,
rapporterar	reports,
norstedt	norstedt,
begått	comitted,committed,
olsson	olsson,
studeras	(is) studied,is studied,
sidan	side,the side,
interstellära	interstellar,
regerande	ruling,
hänvisade	refer,
förblir	remains,remain,
stoft	dust,
träda	fallow,
placerades	placed,
akc	akc,
melankoli	melancholy,
diameter	diameter,
järnmalm	iron ore,
faktiskt	in fact; actually; indeed,
bro	bridge,
läkemedelsverket	medical products agency,
tillsammans	together,
faktiska	actual,
total	total,
absolution	absolution,
stått	stood,
ätten	the dynasty,
debutalbumet	the debut-album,
lämpligt	suitable,
indiana	indiana,
negativt	negative,
supportrar	supports,supporters,
giovanni	giovanni,
fingrar	fingers,
riksväg	national highway,highway,
nku	nku,
lissabonfördraget	treaty of lisbon,lisbon treaty,
kurderna	kurdish,
springer	running,springer,
absorberas	(gets) absorbed,
friheten	freedom; liberty,liberty,
beväpnade	armed,
fascismen	the fascism,fascism,
era	yours,
specialiserade	specialized,
klorofyll	cholophyll,
folkmun	popular lore; popularly,common speech,colloquially,
gloria	gloria,
vackra	beautiful,
ekonomiskt	economic,economical,
sommar	summer,
vers	verse,
indien	india,
felaktigt	incorrect,erronenous,
indier	indians,
enhet	unit,entity,
valborg	valborg,
utlandet	foreign land,abroad,foreign,
gotlands	gotland's,
solen	the sun,sol,
firas	celebrated,celebrate,
firar	celebrates,celebrate,
gillar	likes,enjoy; like,
leonard	leonard,
halland	halland,
sammansatt	composed,
rädd	afraid,
biografer	movie theaters,movie theaters; cinemas,cinemas,
kategorieuropas	category europe,
lag	law,
koreakriget	the korean war,
tjäna	profit,earn,
biografen	the cinema,
orden	the words,
medlemsstat	member state,
vänsterpartiet	leftist party,left-wing party,left wing party,
lämningar	remains,remnants,
massmedia	media,mass media,
dagbladet	daily paper,
över	of,over,
arbetslöshet	unemplyment,
natten	overnight,
office	office,
sovjet	soviet,
exempel	example,for example; for instance; sample(-s),
inspelningarna	recordings,
söderut	south,
blandning	mix,mixture,
japan	japan,
bidra	contribute,
vilken	what,which,
straff	penalty,punishment,
lagets	the team's,
fragment	fragment,
vanligtvis	usually,generally,
band	band,
fredsbevarande	peacekeeping,
bana	course,
they	they,
spelningen	the gig,
bank	bank,
huvudartikel	main article,principal article,
l	l,
dåliga	bad,
diskuteras	discussed,is discucssed,
knutpunkt	hub,
tendens	tendency,
område	area,
carlos	carlos,
germanska	germanic,germanian,
inflytandet	the influence,
koldioxid	co,
voddler	voddler,
däggdjur	mammalian,mammal,
rummet	room,
kejserliga	imperially,
asteroidbältet	the asteroid belt,
därav	thereof,
trafik	traffic,
bruttonationalprodukt	bnp,
oskar	oskar,
vete	wheat,
funktionen	function,the function,
veta	know,
nationalistiska	nationalist,nationalistic,
veto	veto,vetoe,
standard	standard,
förmodligen	probably,presumably,
tillbaka	back,
berör	affect,concerns,
ange	name,
sprit	liqeur,
väldiga	immense,vast,
professionell	professional,
väldigt	very,
förmågan	the ability,
personerna	people; persons,the persons,
föras	taken to,
önskar	wish,
statskupp	coup,
ingmar	ingmar,
synnerligen	remarkably; particularly,particularly,quite,
paret	the couple,
drabbade	suffering,affected,
begränsas	limited,(gets) limited,
begränsar	limits,
ingen	there is no,no,
begränsat	limited,
förklarade	explained,
växthusgaser	greenhouse gas,
inget	no,
john	john,
begränsad	limited,
antisemitismen	antisemitism,anti-semitism,
äter	eat,eats,
militärt	militarily,
albert	albert,
åland	Åland,
kvarvarande	lasting,remaining,residual,
persson	persson,
bojkott	boycott,
kraftverk	power plant,
trupp	troops,troop,
källkod	source,source code,
militära	military,
nedan	below,hereinafter referred to as,
toronto	toronto,
binda	bind,tying,
kronan	kronan,swedish krona,
sonen	the son,
används	use,used,
scenen	the stage,
binds	bound,(is) bound,
byggts	built,
minut	minute,
pelle	pelle,
använda	using,
årens	the year's,
skolorna	the schools,
mannen	the man,
inverkan	impact,influence,
höja	increase,raise,
omvandling	transformation,
framtida	future,
kallades	was called,summoned,
anledningar	reasons,
kalendern	calender,
magnus	magnus,
höjd	height; above,height,
sjukvård	health care,healthcare,
aftonbladet	aftonbladet,the evening paper,
lades	put,
figurerna	figures,characters,
närvaro	attendance,
historisk	historic,historical,
verkar	seems,operates,
maiden	maiden,
bruce	bruce,
utställning	exhibition,
fjädrar	feathers,
verkan	effect,
flygplatsen	the airport,
aminosyra	amino acid,
eviga	eternal,
ägda	owned,
freja	freja,
ägde	tookplace; occured,
bortom	beyond,
läran	teaching,the teaching,
evigt	forever,eternal,
förväxla	mistake,
effekten	the effect,effect,
mitten	middle,mid,
damer	ladies,
lewis	lewis,
hinduiska	hindu,
madeira	madeira,
tilläts	was allowed,were allowed to,allowed,
vintrar	winters,
senare	latterly; later,later,
fortplantning	reproduction,sex,
rankning	ranking,
sättet	manner,way,the way,
 kilometer	kilometer,
sätter	place,puts,sets,
näring	nutrition,
estetiska	aesthetic,
handlar	concerns,
kejsar	emperor,
inställning	attitude,view,
målvakt	goalee,goalkeeper,
variera	vary,
kontinuerlig	continuous,
imperium	empire,
dj	dj,
de	the,
sverigedemokraterna	sweden democrats,swedish democracy,
stalins	stalins,stalin,
watson	watson,
människorna	men,the humans,
orolig	worried,
riktningen	direction,denomination,
du	you,
dr	doctor,dr,doktor,
sattes	was added,
offret	the victim,offering,
runt	around,between,
spridningen	spread,the spread,
konst	art,
splittrades	shattered,split,
offren	victims,
tyngre	heavier,
fågelarter	species of bird,
lasse	lasse,
libanon	lebanon,
kurdiska	kurdish,
vanlig	common,
utförd	completed,performed,
treenigheten	tinity,
förena	combine,unite,
grundarna	founders,
historiens	historys,history's,
präglats	been marked,marked,
utfört	done,
utförs	is done,
sexuell	sexual,
djuret	the animal,
fornnordiska	old nordic,ancient nordic,
fångenskap	captivity,
djuren	the animals,
materialet	the material,
smaken	the flavour,
militärer	soldiers,
we	we,
självständigheten	independance,
intog	seized,
miljö	environment,
jämförelse	comparison,
huvudsakligen	generally,primarily,
militären	the military,
garanterar	ensures,guarantees,
kännetecknas	characterized (by),characterized,
kommer	is,
brad	brad,
gruppens	group (-s),
målningen	milling,the painting,
vecka	week,
graviditeten	the pregnacy,the pregnancy,
kännetecken	distinction,
thierry	thierry,
fångar	prisoners,
tusentals	thousands,
genomför	carry out,
tony	tony,
slaveriet	slavery,
smith	smith,
japans	japans,japan's,
patienten	the patient,
tids	time,
lösning	solution,solution; resolution,
framträdande	apperance,appearance,
hitlers	hitlers,
patienter	patients,
klubblag	club teams,
nära	close,
attacken	the attack,
attacker	attacks,assaults,
fest	festival,party,fest,
juridik	law,
drottningen	the queen,
frekvens	frequency,
bulgariens	bulgaria's,
vagn	wagon,
johansson	johansson,
påstådda	said,alleged,
kupp	kupp,coup (d'etat),
nordöstra	northeast,
klippa	cut,
spanjorerna	the spaniards,spanish,
have	have,
moldavien	moldova,
deltagarna	the participants,participants,
jordbruk	agricultural,
påverkades	was affected by,affected,
själva	self,actual,
våg	road,wave,
patent	patent,
bergskedjor	mountain ranges,
självt	itself,
utgivna	issued,published,
ersattes	was replaced by,replaced,
andelen	share,the share,the proportion,
producerades	was produced,
raid	raid,
hann	reached,managed to (in a period of time),
saddam	saddam,
balkan	balkan,the balkans,
sexualitet	sexuality,
delstater	states,
hand	hand,
delstaten	the state,
hans	his,
bilen	the car,
koncentrerad	concentrated,concentration,
aspekter	aspects,
förlorade	lost,
rörelsen	movement,
kyla	cold,cooling,
riksdag	parliament; diet,parliament,
rör	touch, move(-s),touches,
styrkorna	forces,
mamma	mother,
monaco	monaco,
rörelser	movements,
röd	red,
thc	thc,
gärningsmannen	perpetrator; offender,the offender,culprit,
newton	newton,
kall	cold,
nästan	almost,
kroppens	the body's,the bodies,
goda	good,
enades	agreed,
kalender	calendar,calender,
upptäckte	discovered,
swahili	swahili,swahilli,
världsdel	continent,
så	so,
distributioner	distributions,
påföljande	subsequent,
wright	wright,
havets	sea,
sjunka	descend,
skick	state,condition,
kvinnan	woman,
plasma	plasma,
viking	viking,
förbättra	improve,
föda	give birth; food,give birth,
återgick	returned,returning,
skadorna	injuries,damages,damage,
arab	arab,
fusion	fusion,
indianer	indians,
föds	born,
everton	everton,
engelskans	english,
hepatit	hepatite,hepatitis,heptatitis,
acceptera	accept,
årlig	yearly,
indelning	the subdivision,classification,
indelningen	division,classification,
syfte	view,
samfund	communities,order,
gandhi	gandhi,
transkription	transcript,transcripton,
sixx	sixx,
motsvarighet	equivalent,
korea	korea,
avsätta	unseat,
bort	away,remove,
presidentvalet	presidential elections,presidential election,
borg	tower,
bord	table,
kungar	kings,
humor	humour,
territorierna	territories,
serbiens	serbias,
siffran	number,the number,
vinterkriget	the winter war,
stadsdelarna	districts,neighborhood (-s),
vägar	roads,paths,
bevara	preserve,
fängslades	imprisoned; jailed, gaoled; incarcerated,jailed,
post	not a swedish word,
detta	this,
vunnit	win,won,
upplösning	resolution; dissolution,resolution,
banker	banks,
juryns	the jury's,
jacques	jacques,
återfinns	is rediscovered,
tjänstemän	officals,
lois	lois,
epicentrum	epicentre,
fängslade	inprisoned,confine,
blivande	future,to be,
gemenskapen	the collective,
way	väg,
war	war,
etablerat	established,
hypotes	hypothesis,
skiljas	separate,
motorvägar	highways,motor,
inträffar	occurs,occur,
inträffat	occurred,
partiledare	party leader,
emil	emil,
reser	travels,rise,rises,
studierna	studies,the studies,
finansiering	financiation,
litterär	literary,
långvarig	of long duration,prolonged; lengthy; long,long,
träning	training,practice,
erövra	conquer,
engagerade	dedicated,engaged,committed,
utomlands	abroad,
tesla	tesla,
xiis	xii,
efter	after,
bilderna	the pictures,
xiii	xiii,
moln	cloud,
empati	empathy,
toppen	top,peak,the top,
alltid	always,
möta	meet,
förmåga	abilities,ability,
janukovytj	janukovytj,
knäppupp	knäppup,knäppupp,
arkitekter	architects,
test	test,
götaland	götaland,
konservatism	conservatism,
mött	faced,met,
femton	fifteen,
tottenham	tottenham,
inspelad	recorded,
reglerar	regulates,
regleras	regulated,
rätter	dishes,
hemma	at home,
omgivande	surrounding,surounding,ambient,
rätten	the court,
solens	the sun,
bergmans	bergman's,bergmans,
uppfanns	invented,
tenderar	tend,
datum	date,
nervosa	nervosa,
osäker	insecure,
lider	suffers,
utkämpades	fought,
förhistorisk	prehistorian,
brottet	the crime,the crime; offense; infraction; transgression,
afrikaner	africans,
heller	neither,neither; nor,
rådet	the council,council,
igelkott	hedgehog,
terror	terror,
vänder	turn,
brown	brown,
hannah	hannah,
uttrycka	express,
försörjde	provided,
lättare	easier,
hannar	males,
vegas	vegas,
uttryckt	expressed,
avbröts	canceled,interrupted,
enskilt	individually,
salvador	salvador,
stycken	pieces; parts,
nedsatt	impaired,reduced,decreased; diminished,
datorspel	video game,computer game,
hisingen	hisingen,
levnadsstandard	living standard,standard of living,
frigörs	is released,
ljuset	the light,
ordet	the word,
formella	formal,
litterära	literary,literal,
templet	the temple,temple,
revolution	revolution,
alfa	alpha,
cosa	cosa,
engagerad	engaged,
invandrade	immigrant,
sköttes	operated,handled,
mål	goal,
formellt	formally,formal,
motsatte	opposed,
stimulera	stimulate,
motsatta	opposite,
ungdomar	youths,adolescents,the youth,
tidig	early,
ingick	were included,
kosmiska	the cosmic,
uniform	uniform,
fastigheter	real estates,
utspelar	takes place,set,
versionen	the version,
gener	genes,
oerhörd	tremendous,
marxismen	marxism,the marxism,
kärlek	love,
påstås	claimed,(been) said,allegedly,
påstår	claims,asserts,
genen	gene,the gene,
oerhört	tremendously,
tillträde	access,
antarktiska	antarctic,
sistnämnda	later,
gård	farm,
kemi	chemistry,
avsnitten	the episodes,chapters,
franklin	franklin,
ponny	pony,
istället	instead of,
vinnare	winner,
ekr	ekr,ad,
churchill	churchill,
marken	soil,
extra	extra,
vapnet	the weapon,the weapon; escutheon; coat of arms; arms; badge,
spridit	spread,
ukrainas	ukranian,ukraine's,
förteckning	index,listing,label,
kärnkraftverk	nuclear power plant,nuclear powerplant,
presenterar	presents,present,
upprättade	established,
äktenskapet	marriage,
förkortat	shortened,
territorier	territories,
stabilitet	stability,
regel	rule,
territoriet	territory,
angels	angels,
överhuvudtaget	in general, generally,
fransmännen	the french,french,
parallellt	at the same time,
club	club,
rivalitet	rivality,rivalry,
snabbt	quickly,
enda	only,
målvakten	the goalkeeper,
ämnena	the elements,substances,
närmar	close in,closing,
varför	why,
kolonialismen	the colonialism,colonialism,
feministiska	feminist,
snabba	rapid,fast,
löner	wages and salaries,salaries,
ibm	ibm,
ibn	ibn,
interaktion	the interaction,interaction,
can	can,
erbjuder	offers,
några	a few,
december	december,
nobels	nobel's,
arean	the area,the space,
gentemot	towards,
abort	abortion,
uppstår	occur,
genomgått	experienced,
kritiserar	criticize,
judendomen	the judaism,judaism,
ligan	league,
pojke	boy,
betydelse	significance,
kopplingar	connections,links,
perserna	the persians,persians,
riktlinjer	guidelines,
framgångarna	successes,the successes,
göteborgs	gothenburgs,
gräns	border,
ungern	hungary,hungaria,
förutsättning	prerequisite,
flyttat	moved,
flyttas	is moved,moved,
flyttar	move,
kurt	kurt,
kurs	course,
michel	michel,
ukrainska	ukrainian,
rekordet	the record,
maktens	the power's,
landshövding	county governor,govenror,
ingripa	interfere,
ganska	rather,quite,
ättlingar	descendants,
respektive	respective,
kombination	combination,
generalguvernören	governor-general,governor general,general governor,
fält	field,
skabb	scab,scabies,
utnämndes	was declared,appointed,
därifrån	from there,
bergskedjan	mountain range,the mountain group,
nominerades	was nominated,nominated,
hals	throat,neck,
varav	of which,which,
halt	stop; level,stop,
halv	half,
nog	sufficiently,enough,
författarna	the authors,writers,
komponenter	components,
begränsa	limit,
jorden	the earth,earth; earth; underground,
nou	nou,
rakt	straight,
now	now,
dödsstraffet	capital punishment; death penalty,the death penalty,
hall	hall,
frihet	freedom,
james	james,
språk	language,
främmande	foreign; alien,foreign,
antyder	indicates,
stockholm	stockholm,
januari	january,
drog	draw,pulled,
aspergers	downs syndrome,aspergers,
em	european championship,
sektorn	the sector,
citat	quote,
ej	not,no,
ed	ed,
eg	ec,
utbrett	wide,widespread,
spåra	track,trace,
strålningen	the radiation,radiation,
ex	ex,
kroatiska	croatian,
et	et,
kant	kant,edge,
fuglesang	fuglesang,
ep	ep,
premiärministern	the prime minister,
er	you,
album	album,
teorier	theories,
återkommande	recurring,
videon	the video,
hustrun	the wife,
kortare	shorter,
stallone	stallone,
hellre	rather,
koffein	caffein,
genetisk	genetic,
taget	a time (practically; virtually; any; at all),
marino	marino,
marina	marine,
betraktades	considered,regarded,
british	british,
domen	verdict; judgement,
allmänheten	public,general public,
arbetsgivare	employers,
blind	blind,bank,
xi	xi,
förändrats	changed,
derivatan	the derivative,
ring	ring,
bergqvist	bergqvist,
våglängder	wavelengths,wave lengths,
omtvistat	contentious,disputed,controversial,
priser	prizes,
national	national,
sheen	sheen,
dessutom	furthermore; moreover, additionally; likewise,furthermore,
satsningar	investments,resources,
färre	fewer,less,
spelningar	tour,gigs,
nödvändig	necessary,essential,
fascisterna	the fascists,the facists,
delats	been awarded,
television	television,
europeisk	european,
sidorna	the pages,pages,
utbyggda	expanded,expand,
ändrades	changed,
grundad	founded,
craig	craig,
statsminister	prime minister,
faktor	factor,
kairo	cairo,
grundat	founded,(was) found,
grundar	bases,based,
grundas	is based,based,
anger	gives,
anges	mention,specified,
hjälp	help,
hör	belong,
skär	skerry,
fortsatta	continued,
etiopiska	ethiopian,
bönor	beans,
hög	high,
skäl	reasons,reason,
kategoriorter	category visited,
numera	now,nowadays,
successivt	successively,progressively,
bön	prayer,
bekostnad	expense,
dvärgar	dwarves,dwarfs,
glödlampor	lightbulbs,light bulbs,
användning	use,use; usage,
america	america,
på	on,in, on, at,
lyfter	lifts,lifting,
norrmän	norwegians,
nordligaste	northermost,northern,northernmost,
parlamentets	the parliament's,
runda	round,
orsaka	cause,
abraham	abraham,
skapats	was created,
doktor	doctor,
kyrkorna	the churches,
nazisternas	the nazi's,
enighet	unity,
colombo	colombo,
teori	theory,
perfekt	perfect,
mannens	man's,
rötter	roots,
varmblod	warmblood,warm-blooded,
adolf	adolf,
billiga	cheap,
huskvarna	huskvarna,
epoken	the epoch,
dagbok	diary,
sierra	sierra,
mörk	dark,
sydligaste	southernmost,most southern,
uppståndelse	resurrection,
tornet	the tower,
riddare	knight,
samuel	samuel,
mission	mission,
ambitioner	ambitions,
folkomröstning	referendum,
marxistisk	marxist,marxistic,
tävla	compete,
handlingar	actions,
drabbas	suffer,troubled with,
facupen	fa cup,fa-cup,
tvingade	forced,
bushadministrationen	the bushadministration,bush administration,
länge	long,
storstäder	metropolises,
osbourne	osbourne,
övergången	the transition,transformation,
sport	athletics,sport,
långsammare	slower,
depressionen	the depression,
konstaterade	concluded,established,stated,
ladin	ladin,
depressioner	depressions,
israels	israel's,
import	import,
kommunismens	the communisms,the communism's,
katastrofen	catastrophy,the catastrophy,disaster,
sträcka	distance,
ronja	ronja,
ordspråk	saying,
flygande	flying,
männen	the men,men,
utgivningen	release,the publication,the release,
verket	plant; indeed,plant,
hendrix	hendrix,
verken	wroks,
utgavs	was published,
samtal	conersation,
monicas	monica's,
representativ	representative,
bördiga	fertile,
placerad	placed,
smålands	smaland's,
kristinas	kristina's,
feminismen	feminism,
ståndpunkt	standpoint,
nils	nils,
comet	comet,
placerar	place,places,
placeras	placed,
utnyttja	use,
avskaffande	abolition,abolishment,
dömande	sentencing,judging,
lägenhet	appartment,
bomull	cotton,
riksrådet	privy council; council of state; crown council; senate,
östtyska	east german,
överlever	survives,
handlande	action,
långfilm	feature film,
oliver	olives,
välstånd	prosperity,
sättas	turn,
karlstads	karlstad's,
sker	happens,
oden	oden,
knappt	barely,
socialdemokrater	social democrats,
dräkt	costume,outfit,
observera	note,observe,
utförda	made,
riktningar	directions,direction (-s),
elvis	elvis,
funnits	been,
anslöt	joined,
ytan	the area,
uefacupen	the uefa champions league,uefa europa league,
rapporter	reports,
prinsessan	the princess,princess,
rapporten	the report,
polens	polands,
ordningen	the order,
ändå	still,
ansikte	face,
tjeckien	czech republic,the czech republic,
eran	era,
beläget	located,
inslag	elements,
finanskrisen	the financial crisis,
tänkande	thinking,
behandlade	was treated,
kvarter	block,
kenya	kenya,
västerländska	western,
katalanska	catalan,
helium	helium,
grundade	founded,based,
infödda	natives,
slaget	the strike,
långt	far,
orsakade	caused,
programvara	software,
media	media,
långa	long,
talmannen	speaker of the riksdag,
homosexualitet	homosexuality,homosexuallity,
kromosom	chromosome,
pesten	the plague,death,
lite	little,
speciella	special,
offensiven	offensive,the offensive,
begär	requests,
skivbolaget	record label,the record company,
acdc	ac/dc,
omfattande	wide-ranging,large,massive; extensive,
målningar	paintings,
omfattas	comprise,
speciellt	particularly,
omgående	immediate,
ekonomisk	economic,
tradition	tradition,
fredspris	peace prize,
skånes	scania's,
erkänd	acknowledged,
erkänt	recognized,
flaggor	flags,
mynning	outfall,muzzle,mouth,
forskarna	the scientists,
skandinaviska	scandinavic,scandinavian,
tydlig	clear,obvious,
framgången	the success,
eleverna	the pupils,the students,
lagerkvist	lagerkvist,
spänningar	tensions,
nazismen	nazism,
euron	the euro,
lade	laid,seized,
ditt	your,
strävar	striving; aiming (to; for),strives,
irland	ireland,
arbeta	work,
passiv	passive,
stund	while,
östergötland	Östergötland,
selma	selma,
amy	amy,
rebecca	rebecca,
symbolisk	symbolic,
strävan	will,the quest,endeavor,
skilda	seperated,separate,
miniatyr|en	a minature,
skilde	divided,there was a separation,
varandra	each other,
nationellt	nationally,
t	t,
låga	low,
eddie	eddie,
lågt	low,
präglades	imprinted,marked,
stånd	in the context: (make) the war happen,position,
fönster	window,
slår	states,beats,
användbara	usable,useful,
sålts	sold,
indikerar	indicates,
frigörelse	liberation,
berodde	depended,depended upon,
agera	act,
strindberg	strindberg,
utskott	committee,organ,
bestämt	decided,
nsdap	nsdap,
inuti	inside,
växa	grow,
kategoriledamöter	category: members,
bestäms	is decided,
kaffet	the coffee,
francis	francis,
övertygad	confident,
ideologi	ideology,
central	central,
bidraget	contribution,
sri	sri,
kompositörer	composers,compositors,
torget	square,the square,
bidragen	the contributions,contributions,
efterkrigstiden	the post-war period,post-war era,
kapten	captain,
klassiker	classic,
utbildade	educated,
karriär	career,
area	area,
satsade	bet,
sats	theorem,
stark	strong,
start	start,
anställd	employed,hired,
danska	danish,
specifika	specific,
likväl	nevertheless,still,as well,
gånger	times,
fastställa	determine,confirm,
hawking	hawking,
tunisien	tunisia,
guillou	guillou,
wailers	wailers,
sämsta	worst,
gången	time,
traditionerna	traditions,the traditions,
expeditionen	the expidition,
spänner	span,
minne	memory,
engelskan	the english,
indelningar	divisions,classifications,
minns	remembers,remember,
miguel	miguel,
bilmärke	car make,make of car,
expeditioner	expeditions,
kostar	costs,
kungen	the king,
grammis	grammy,
sveriges	swedens,
godkände	approved,
styrde	steered,
knut	knut,knot,
transportera	transport,
nere	down,
drycker	beverages,
efteråt	afterwards,
upphovsman	author,
köper	making,
knä	knee,
drift	drift,
översätts	translate,is translated,
massachusetts	massachusetts,massachussetts,
röda	red,
bandmedlemmarna	band members,have,
skuggan	shadow,the shadow,
tjänare	servant,
handelsmän	merchants,
morgonen	the morning,
färdas	travels,
susan	susan,
olympiastadion	olympa stadium,olympic stadium,
eriksson	eriksson,
beskrivningar	descriptions,
bäst	best,
messi	messi,
öknen	the desert,
loppet	the race,
antoinette	antoinette,
griffin	griffin,
armar	arms,
lämpliga	suitable,
påbörjades	commenced; begun,initiated,was started,
foster	fetus,
fästning	fortress,
skiljer	differs,is different; differ,different,
kolonierna	colonies,
får	can,allow,
verk	work,works,
osv	etc.,
tredje	third,
heaven	heaven,
sverige	sweden,
behöver	need,
louis	louis,
mild	mild,
industrialiseringen	indutrialization,industrialization,
resan	the trip,
rasism	racism,
magdalena	magdalena,
skiva	record,disc,
fåglarnas	the birds',birds,
egendom	property,
kritiserats	criticized,critized,
bestämde	determined,chose,
orgasm	orgasm,
markerade	marked,
trupper	troops,
utåt	outwardly,out,
pythagoras	pythagoras,
tvskådespelare	tv actor,
besöker	visit,visits,
bedrev	managed,
fjärde	fourth,
förbjuden	smoking,
bernhard	bernhard,
förbjuder	forbids,
misstänkta	suspected,
inblandad	mixed,
klassificera	classifying,
irak	iraq,
ersatt	replaced,
iran	iran,
genomförde	carried out,
ersättare	replacement,
kronor	kronor,
observeras	observed,is noticed,is observed,
uttalat	outspoken,expressed,
lämna	leave,
uttalas	be pronounced,
arena	arena,
medarbetare	coworker,
vår	spring,
krigen	the wars,wars,
stulna	stolen,
minst	at least,
boxning	boxing,boxing; pugilism,
sagor	fairytales,tales,fairy tales,
kriget	the war,
hoppades	hoped,
perspektiv	perspective,
då	then,
globen	the globe,
nazityskland	nazi germany,
gick	went,passed,
grunda	found,
dalarna	dalarna,
ökat	increased,
nukleotider	nucleotides,nucleotide,
familj	family,
avsedd	intended,
simba	simba,
arrangemang	arrangement,
taket	the roof,
tillät	allowed,
etablerad	established,
förlängningen	elongation,
planen	the field,the plan,
bolagets	company's,the corporation's,
representeras	represented,
representerar	represents,
massan	mass,
kurdistan	kurdistan,
reptiler	reptiles,
okänt	unknown,
utökat	extended,
blodtryck	blood pressure,
ständiga	permanent,constant,
latinamerikanska	latin-american,latin american,
räknat	calculated,counted,
räknar	counts,counter,
räknas	counted,are counted,
lagstiftande	legislative,legislating,legislation,
ständigt	always,constant,
nina	nina,
företeelser	phenomena,
gazaremsan	gaza strip,the gaza strip,
ombord	onboard,
livslängd	life expectancy,
fronten	front,the front,
rapporterade	reported,
kejsardömet	empire,
partner	partner,
fatta	make,
herrens	lord,
zanzibar	zanzibar,
serber	serbs,
ledger	ledger,
linköping	linköping,
smitta	infection,
reidars	reidars,reidar's,
kung	king,
samarbetet	cooperation,the collaboration,
utför	perform,
turkarna	the turks,
torde	could,should,
fastän	although,
försök	expirements,
fd	ex,
ff	ff,
invasion	invasion,
samarbeten	cooperations,collaborations,
fn	un,the un,
stabil	stable,
vattenkraft	water power,hydroelectric power,
kostnaden	cost,
byggandet	the building,
skivan	record,the record,
enzymer	enzymes,
allmänna	general,
kognitiv	cognitive,
segrar	wins,victories,
skiljs	separated,separate,
kostnader	costs,expenses,
dream	dream,
nämnts	mentioned,
tillgångar	assets,
helt	totally,
helgdagar	holidays,
tornen	towers,
hela	entire,
maffian	mafia,
hell	hell,
kombinerade	combined,
eros	eros,
hundratusentals	hundreds of thousands of,hundreds of thousands,
romance	romance,
kusterna	the coasts,
antagits	adopted,
systems	systems,
österrikes	austria's,austrias,
mahatma	mahatma,
musikalisk	musical,
bytte	changed it's,swapped,
elden	the fire,
lyckas	succeed,
konstitutionella	constitutional,
greps	was arrested,(was) arrested,
dyrt	a high price,expensive,dearly,
petter	petter,
närmare	close to,
fullt	full; fully; completely,completely,full,
fulla	full,complete,
skrivit	written,wrote,
strålning	radiation,
kontinentens	the continents,
ifk	ifk,
etnisk	ethnic,
positionen	the position,
positioner	positions,
rättvisa	justice,
försäljning	sales,sale,
aktörer	players,actors,
robert	robert,
bodde	lived,
lungorna	the lungs,
stödet	support,the support,
stöder	supporting,supports,
känna	know,
efternamn	last name,lastname,surname,
utredningen	the investigation,
heroin	heroine,
känns	feels,
delningen	division,pitch,
vasas	vasas,vasa's,
svarade	answered,accounted (for); answered,
etnicitet	ethnic,
skogen	forest,
skilja	seperate,differ; differentiate,separate,
förbättrade	improve,
underhåll	support,allowance,
ytterligare	further,additional,
sänder	broadcast,transmits,
sändes	was sent,
utvecklats	developed,
synen	the view,sight,
etiska	ehtical,
arsenal	arsenal,
minoritetsspråk	minority language,minority,
fabriker	plants,factories,
helsingborgs	helsingborg's,
taggar	spikes,thorn, twig,
synes	appears,
miss	miss,
rygg	backs,back,
deltagare	contestant,participiant,
kanada	canada,
kongresspartiet	congress party,indian national congress,
station	station,
parlamentsvalet	parliament election,election to parliament,
nigeria	nigeria,
brittiska	british,
luminositet	luminosity,
nominerad	nominate,nominated,
åkte	went,relegated,
förnuftet	the common sense,
brittiskt	brittish,british,
tvungen	forced,forced (to),
bildande	formation,founding,
växterna	plants,
brasiliens	brazil's,
långsamt	slowly,
einsteins	einsteins,
andersson	andersson,
värden	values,
värdet	the value,
signifikant	significant,
gren	branch,
familjerna	families,
öde	fate,
avancerade	advanced,
charlotte	charlotte,
bestämdes	was decided,decided,was determined,
teslas	tesla's,
genomgripande	good,comprehensive; radical,
medeltemperaturen	median temperature,
tvärtom	on the contrary,contrary to,
brittiske	british,
militär	military,
demokratin	the democracy,
vädret	the weather,
liberalismen	the liberalism,
lik	similar,alike,
liv	life,
ledde	resulted,led,
herre	lord,master; lord,
avseenden	respects,regard,
jämföras	compared,
mexiko	mexico,
logotyp	logotype,
säsongens	the seasons,
bistånd	aid,
kap	chapter,cape,
kongress	congress,
utgör	make up,constitutes,
himlakroppar	celestial bodies,
kokain	cocaine,cocain,
polacker	polish,poles,
klädd	clothed,
räknade	counted,
recensioner	reviews,
rådde	prevailed,was,
två	two,
osäkra	insecure,uncertain,
ingenting	nothing,
jupiters	jupiter's,
möjligen	possibly,
muslimsk	muslim,muslim; muslem,
integritet	integrity,
justice	justice,
humanistiska	humane,humanistic,
åländska	Åland swedish,
ikon	icon,
lönneberga	lönneberga,lonneberga,
darwin	darwin,
ingå	be a part,be included in,
dominans	dominant,dominance,
arabvärlden	the arab world,
tillhört	belonged,
utrikes	foreign,
tillhöra	belong to,
alexander	alexander,
restauranger	restaurant,restaurants,
avsaknaden	absence,
dömdes	sentenced,was convicted,
vilket	which,
målare	painter,
tolkiens	tolkien's,
västkusten	the west coast,west coast,
grunden	basis,
allmänt	generally; public,commonly,
maurice	maurice,
bakgrund	background,
tidigare	earlier,
ändamål	purpose,
mörkare	darker,
flyter	flows,
gravitation	gravitation,
haddock	haddock,
upphovsrätten	copyright,
pjäser	plays,
löst	solved,1st sentence: loosely; 2nd & 3rd: solved,
produkten	the result,product,
chansen	chance,
allvar	earnest,
likhet	similar,resemblance,like,
utsträckning	extent,
köket	the kitchen,
revolutionen	the revolution,revolution,
länk	link,
produkter	products,
lejonet	the lion,
anor	lineage; ancestry,
viljan	will,
slavar	slaves,
kyrkliga	religious,
bott	lived in,
läsaren	the reader,reader,
uppfylla	satisfy,fulfill,meet (requirements),
betydde	meant,ment,
derivata	derivative,
scientologikyrkan	church of scientology,
sokrates	sokrates,socrates,
vintertid	winter-time,
händerna	hands,
merparten	most,the majority,larger part,
minskade	was reduced,
enheten	the unit,
enheter	units,
kuster	coasts,
konsensus	consensus,
gestalt	character,figure,
walter	walter,
isolerade	isolated,
handlingen	the plot,the story,
budgeten	the budget,
anthony	anthony,
livet	the life,life,
delades	shared,divided,split,
genomförs	implemented, carried through,conducted,
socialism	socialism,
belgrad	belgrade,
hegel	hegel,
läser	are reading,
diktator	dictator,
mängden	amount,the amount,
tillfället	to the case,
slutar	ends,end,
slutat	ended,
uttryckte	expressed,
nationalitet	nationality,
klippiga	rocky,
sorter	kinds,types,
bärande	wearing,leading,fundamental; wearing; supportive,
lagar	laws,
tillfällen	oppertunities,jobs,
kombineras	combined,
staffan	staffan,
kombinerat	combined,
ändra	change,
deltagande	participation,
sammanlagt	a total of,
nöd	distress,
kombinerad	combined,
inledde	started,
folkslag	kind of people,
kungahuset	royal house,
bon	bon,
anklagats	accused,
 km	kilometers,
kommunicera	communicate,
förlag	magazine,
chris	chris,
seglade	sailed,
armenien	armenien,armenian,
svealand	svealand,
bob	bob,
kurdisk	kurdish,
stjärnorna	stars,
präglas	characterised,characterized,
flygplan	aircraft,airplane,
nutid	present day,present,
präglad	characterize,marked,characterized,
innersta	innermost,
feminister	feminists,
departement	department,
njurarna	the kidneys,
tortyr	torture,
skal	shell,
fredliga	peacefull,peaceful,
inlett	started,ushered in,
uppfinnare	inventor,
kallblod	cold blood,draught horse,
taiwan	taiwan,
henne	her,
gänget	the group,the gang,
nikki	nikki,
välkända	well known,
varuhus	warehouse,
egenskap	trait,ability,seeks,
djup	deep,
marco	marco,
bestå	exist,
återställa	restore,
lika	similar,alike,equal,
gör	does,makes,
kulturen	the culture,
enklare	easier,simpler,
kulturer	cultures,
gitarristen	the guitarist,guitarists,
unga	young,
immigranter	immigrants,
innan	before,
uppvärmningen	the warmup,heating,the warm-up,
releasedatum	release date,
dylikt	such,
koden	the code,
infektion	infection,
criss	criss,
gandhis	gandhi's,
terminologi	terminology,
unge	young,kid,
donna	donna,
mycket	very,much,
kommenterade	commented,
byggnader	buildings,structures,
biträdande	assisting,
våldet	the violence,violence,
economic	economic,
byggnaden	building,the building,
syndrom	syndrom,
sammanhängande	continous,connective,
skapat	created,
världsarvslista	world heritage list,
vilda	wild,
skapar	creates,
skapas	creates,
faktorn	factor,
enormt	gigantic,
bägge	both,
kejsarens	the emperor's,emperors,
run	run,
steg	step,
rum	(took) place,
sten	stone,
mellankrigstiden	interwar years,time between the wars,interwar period,
stjärnans	star's,the star's,the stars,
offside	offside,
freddie	freddie,
führer	fuhrer,fuehrer,
förtroende	confidence,trust,
myndighet	authoroty,authority,
övergick	transended,went over,
linjen	the line,
etablerade	established,
fysiologiska	physiological,
efterträdare	successor,
refererar	refer (to),references,
linjer	routes,lines,
edvard	edvard,edward,
länderna	the countries,
ändringar	edit,starts to process,changes,
ida	ida,
fåtal	few,a few,
stanna	stop,stay,
egenskaper	characteristics,charactiristics,qualities,
ön	the island,
öl	beer,
reaktorer	reactors,
institut	institution,
emellan	inbetween; between,between,
överst	at the top; uppermost,
föreningen	association,the association,
fokuserade	focused,
ligga	lies, lie,lie,
spänningen	voltage,
visas	is showed,shown,
visat	shown,
heritage	heritage,
spridd	widespread,spread,
jonsson	jonsson,
ledamot	member,representative,
strukturen	the structure,
japanerna	japanese,
spektrumet	spectrum,
larry	larry,
strukturer	structures,
drabbats	affected,afflicted,
skådespelaren	actor,
skull	sake,
ute	out,
nyval	re-election,new election,
skuld	debt,guilt,
malin	malin,
trafikerade	traffic,frequent,
  km²	square kilometre,km2,
politik	politics,
förbjöds	forbidden,
chelsea	chelsea,
ligacupen	league cup,
monarki	monarchy,
ihåg	remember,
avsåg	meant,intended,mean,
voltaires	voltaire,
sydkorea	south korea,
hårdrock	hard rock,hardrock,
igenom	through,
krigets	the war's,war,
sjunde	seventh,
musikens	the music's,
berättat	told,
relationerna	the relationships,relations,
berättar	tells,
berättas	(as) told,told,
korn	korn,barley,grains,
rester	remains,residues,
dras	draw,make (assumptions, references),
drar	earn,
framstående	prominent,
william	william,
drag	trait; characteristic; feature,move,characteristic,
mästare	master,
matematiska	mathematical,
resten	the rest,
vindar	winds,
kors	cross,
närmaste	closest,
samarbetade	collaboration,
enade	united,
medför	entails,result,
dvd	dvd,
officerare	officer,
tunga	heavy,tongue,
heath	heath,
tillfälliga	temporary,
folkliga	popular,
svt	svt,
dvs	(det vill säga) namely that,
skyskrapor	high rise buildings; sky scrapers,
bonniers	bonnier's,bonniers,
höst	autumn,
placera	position,place,
indiska	indian,
katt	cat,
företeelse	experience; phenomenon; feature,phenomenon,
ge	give,
tänker	thinking,
go	go,
träd	tree,
kate	kate,
världsrekord	world record,
baron	baron,
uppgörelse	agreement,deal,
tillhör	belongs,
flitigt	actively,
dröjde	slow,was not until,not until,
sålt	sold,
ännu	still,yet,
rinner	running,flow,
kommunismen	communism,
försvarsminister	minister of defence,
michael	michael,
ryan	ryan,
utbredning	distribution,distrubution,
tidszoner	time zones,
jönköping	jönköping,
stift	diocese,
akut	urgent,acute,
socialdemokratiska	social democratic,
öresund	the sound,
derivator	derivative,derivatives,
mussolinis	mussolini's,
honan	the female,female,
geologiska	geological,
visserligen	certainly,
direkta	direct,
intervjuer	interviews,
börjar	starts,starts to,
börjat	started,begun to,begun,
geologiskt	geological,
svagare	weaker,
kinas	china's,chinas,
erövringar	conquests,
hansson	hansson,
bjöd	invited,
polen	poland,pole,
byttes	changed,was exchanged,
genombrott	breakthrough,
cell	cell,
experiment	experiment,
förhistoria	prehistory,
valen	the elections,
gamla	ancient,
utrikespolitiken	the foreign policy,
gamle	old,
offentlig	public,
innerstaden	inner city,
orsaker	causes,
gåva	gift,
eminem	eminem,
uppgick	total,
ryska	russian,
händelser	happenings,
innebandy	floorball,
västerut	westward; west,westwards,
chans	chance,chanse,
överlevnad	survival,
förening	union,
dopamin	dopamine,
uppfinningar	inventions,
avsedda	aimed,intended,
färöarna	the faroe islands,
vuxen	adult,
italienska	italian,
genetiska	genetic,
personen	the person,
utdöda	extinct,
genetiskt	genetically,genetic,
kunde	could,
stärka	strengthen; bolster,
oktober	october,
sjunger	sings,singing,
starten	the start,
about	about,
invigningen	the opening,
huxley	huxley,
misslyckades	failed,
släppte	released,
debutalbum	debut album,
microsoft	microsoft,
släppts	released,
mottagaren	the receiver,the recipient,
guds	god's,
kenny	kenny,
planerade	planned,
halloween	halloween,
beslöt	decided,
studioalbum	studio album,
talat	spoken,spoke,
fördelningen	distribution,
talas	spoken,
talar	speaks,speak,
romantikens	the romanticism,
tåget	the train,
georg	georg,
tågen	the trains,
sovjetunionen	the soviet union,soviet union,
fälttåg	crusade,campaign,
ferdinand	ferdinand,
folkmängd	population size,population,
kronprinsen	crown prince,the crown prince,
oroligheter	unrest,
fara	danger,
uttalet	the pronounciation,
svenskar	swedish,
dödlig	mortal,
fart	speed,
fars	father's,
utfördes	carried out,preformed,
ringde	called,
österrikiska	austrian,
säljer	sells,
reagerar	reacts,
gått	gone,
encyclopedia	encyclopedia,
förstärka	strengthen,
kungliga	royal,
kapital	capital,
obelix	obelix,
fungerade	working,
presidenter	presidents,president,
offentliga	public,
förstördes	was destroyed,
någonting	anything,
presidenten	the president,
offentligt	public,publicly,
öarna	the islands,
verklighet	reality,
belopp	amounts,
monarken	the monarch,monarch,
begick	commited,committed,
kyrkor	churches,
insekter	insects,
allting	everything,
filosofiska	philosophical,
naturgas	natural gas,
konserten	the concert,concert,
zagreb	capital of croatia,zagreb,
ägna	spend,devote,
läror	teachings,
front	front,
konserter	conserts,concerts,
dikt	poem,
intäkterna	the revenues,proceeds,the revenue,
miniatyr|px|den	miniature,
hunden	the dog,
kläder	clothes,
räckte	enough,
finnas	(be) found,exists,
mode	fashion,
förmågor	abilites,abilities,
täcker	covers,
stadsparken	city park,stadsparken,
föreslogs	proposed,
illuminati	illuminati,
flyg	airforce,air,
skolgång	school attendance,
 procent	percent,
stiger	rises,
skov	forestry,episode,relapse,
skor	shoes,
uppfattar	sees,percieves,interpret,
flyr	flees,escapes,
entertainment	entertainment,
förutom	besides; in addition to; aside from,
islamisk	islamic,
deltagit	participated,
samarbetat	collaborated,
max	max,
solsystem	solar system,
vinter	winter,
omfatta	cover,
torres	torres,
frånträde	relinquishment,withdrawal,
bilder	pictures,
lycka	happiness,
lida	suffer,
bilden	the image,
förstod	understood,
förbund	union,league; alliance; union; compact; covenant,
kommunala	municipal,
florida	florida,
banor	line,
benämnas	named,entitle,
strida	fight,
tillgången	access,
tigrar	tigers,
partierna	political parties,
riksdagsvalet	parliamentary election,election to parliament,
ursprungsbefolkningen	the native population,indigenous population,
minoritet	minority,
brandenburg	brandenburg,
för	to; for,for,
peters	peters,
undervisade	taught,
spaniens	spain's,
boken	paper,the book,
mao	mao,
kulturarv	culture heritage,cultureheritage,cultural heritage,
final	final,finite, final,
zeeland	zeeland,
nilsson	nilsson,
belgiska	belgian,
hasch	hashish,
emellertid	however,
styrelseskick	form of government,
lista	list,
definierat	defined,
definieras	defined,is defined,defines,
definierar	defines,
arbetade	worked,
inbördes	intermutual,
israelisk	israeli,
ber	ask,asks,
bet	bit,
julian	julian,
hjärna	brain,
bordet	the table,desktop,
varade	lasted,
tredjedelar	thirds,
visor	songs,
förlorades	was lost,
släkt	pettigree,family,
attackerna	attacks,the attacks,
runorna	the runes,
röst	voice,
förblev	remained,
jorge	jorge,
galleri	gallery,
regn	rain,
montana	montana,
kvarstår	remains,
regi	direction,
tyskar	germans,
sändas	broadcast,
nå	reach,
överföring	transfer,
skogar	forests,
långtgående	far-reaching,
platon	platon,
parker	parker,
fiktiv	fictive,
tolkien	tolkien,
fynden	finds; findings,
församling	congregation,
passa	take the opportunity,fit,
parken	park,the park,
hade	had,
basen	the base,
radioaktivt	radioactive,
baser	bases,
gemensam	joint,common,
härskare	ruler,
förbli	remain,
varit	has been,been,
partnern	partner,the partner,
aspekt	aspect,
psykologin	the psyhology,
boris	boris,
klassiska	classic,
förespråkare	spokesman,
inbördeskrig	civil war,
omloppsbana	orbit,
michigan	michigan,
området	the area,
inflytelserika	influential,
klassiskt	classical,classic,
häst	horse,
områden	areas,
städerna	the towns,
karriären	the career,
älskade	loved,loved; beloved,
gray	gray,
evolution	evolution,
processer	processes,
tillgång	access,
grav	grave,
influensa	influenza,flue,
också	also,
grad	grade,
kvadratkilometer	square kilometer,square kilometers,
processen	process,the process,
vänt	turned,
sydafrika	south africa,
västindien	west india,
förband	units; formations; bound (themselves),
neutralt	neutral,
landsting	county council,
stats	state's,
tenn	tin,
individens	individual's,the individual's,
flicka	girl,
gotiska	gothic,
staty	statue,
state	state,
företagets	the company's,the corporation's,
ken	ken,
högra	right,
ersätta	replace,
sovjetiska	soviet,sovjet,
benämningen	the designation,the name,label,
merry	merry,
jobba	work,
befälet	the command,command,
problem	problem,
tjänster	services,
kaffe	coffee,
odens	odin's,oden's,
vulkaner	volcanos,volcanoes,
framgångsrika	successful,successes,succesful,
trädde	come into effect,entered,
varierade	varied,
älskar	loves,
stratton	stratton,
framgångsrikt	successful,successfully,
partiklar	particles,
jersey	jersey,
uppsättning	equipment,
fördelar	advantages,share,
fördelas	be allocated,distribute,
torn	tower,
kategoribrittiska	category: british,
leipzig	leipzig,liepzig,
johans	johan's,
genre	genre,
johann	john,
kings	king's,
sammanhang	context,
christer	chris,christer,
liberala	liberal,
trycket	pressure,
sara	sara,
fokusera	focus,
äldre	older,
poet	poet,
påminde	reminded,
poes	poe's,poes,
pontus	pontus,
vinci	vinci,
affärer	business,
spanska	spanish,
spaniel	spaniel,
spanien	spain,
humör	temper,mood,
strömningar	tendencies,sentiments,
kanarieöarna	canary islands,the canary islands,
 meter	metre,meter,
erbjuda	offer,
könsorganen	sex organs,the reproductive organs,
utgjorde	made up,comprised; consisted of,
platons	platon's,platos,
reaktion	reaction,reaction reaction,
nordens	the scandinavian countries',nordic,
rysslands	russia's,
enkel	simple,plain,
erkänner	admits,
feber	fever,
demo	demo,
rättigheter	rights,
mysterium	mystery,
nordirland	north ireland,
måleri	painting,
alfabetisk	alphabetical,
revir	turf,territory,
reformationen	the reformation,
parti	party,
friidrott	track and field,
autism	autism,
varmed	whereby,
begav	went,went (to),traveled,
griffon	griffon,
förebyggande	preventing,preventive,prevention,
korrekta	correct,
flygbolag	airline,
anka	anka,duck,
nationens	the nation's,
rankas	ranks,rank,
införa	introduce,
eklund	eklund,
nämligen	namely,
infört	introduced,
alperna	the alps,
lagring	storage,
flickan	girl,the girl,
strömmen	the stream,
grenar	branches,
i	in,
kärleken	the love,
theodor	theodor,
europarådet	council of europe,european council,
onda	evil,
rösta	vote,
störta	rush,crash,
sänds	sends,
sofia	sofia,
omkom	perished,died; was killed,
sofie	sofie,
förekommer	occurs,
sända	broadcast,send,
sände	sent,
vida	wide,
jeff	jeff,
särskilt	particulary,especially,
natt	night,
nato	nato,
sweet	söt,
titta	watch,look,
bebyggelsen	building,human settlement,settlement,
katolska	catholic,
utan	without,
sanning	truth,
vanligare	more common,
historia	history,
definitivt	unavoidable,definitely,
historik	history,
klassificering	classification,
använts	was used,
lincoln	lincoln,
norges	norway's,
fernando	fernando,
martin	martin,
page	page,
regeringar	governments,
lager	layer,
nationalpark	national park,
vardagliga	ordinary,
pojkarna	boys,the boys,
förlusterna	the losses,
vardagligt	everyday,
förenklat	simplified,made easier,
omöjligt	impossible,
skorpan	crust,
peter	peter,
lagen	the law,law,
moskva	moscow,
skrifter	writings,
 km²	kilometres,
kaspiska	caspian,
hyser	has,accomodates,holds,
folkets	the people's,
alliansen	the alliance,
förde	led,
skriften	writings,
ledd	led,
hinder	obstacle,
motsättningar	contradictions,oppositions,frictions; clashes,
meddelade	informed; announced,stated,
samlades	collected,gathered,were united,
journal	journal,
reza	reza,
kromosomer	chromosomes,
halvön	the peninsula,
usas	usa:s,
keramik	ceramic,ceramics,
föremål	subject,
beslutade	decided,
samlats	gathered; collected,
göteborg	gothenburg,
polisens	the police's,
troligen	probably,likely,
synsätt	effects,viewpoint,
hävdade	claimed,
mytologi	mythology,
betydelsefulla	significant,
glenn	glenn,
washington	washington,
räddade	saved,
tendenser	tendencies,
längsta	longest,
hammarby	hammarby,
museum	museum,
djävulen	the devil,
realiteten	reality,
afrika	africa,
oändligt	infinitely,
distinkt	distinct,distinctive,
cricket	cricket,
står	standing,star,
instiftade	established,created,
neutral	neutral,
ho	ho,
behov	necessary,
hc	h.c.,h.c,
ha	have,
samtida	contemporary,
avled	deceased,
svarta	black,
stål	steel,
fysik	physics,
allierad	allied,
dator	computer,
pippin	pippin pippin pippin,pippin,
komiker	comic,comedian,
förslaget	proposition,the suggestion,
hästar	horses,
invandring	immigration,
bitar	bit,pieces,
farlig	dangerous,
ordbok	glossary,dictionary,
erik	erik,
själ	soul,
motsvarar	comparable,corresponds to the,
eric	eric,
diego	diego,
omväxlande	varied,
sänktes	sunk,
moderaterna	the moderate,the moderates,moderates,
speciell	special,
mineraler	minerals,
hotade	threatened,
vulkaniska	vulcanic,
enastående	exceptional,
stat	state,
revolutionära	revolutionary,
stad	city,
musikvideon	music video,
resulterade	resulted,
stan	town,
ockupationen	the occupation,
hjärnan	brain,the brain,
stam	strain,tribe,
etiken	the ethic,ethics,
förekomma	occur,be found,
inser	recognize,realizes,
klass	grade; class,
alkohol	alcohol,
blogg	blog,
konsumtion	consumption,
hinner	reach it (in time),have time to,
felaktig	incorrect,false,
auktoritära	authoritarian,
andra	other,
nyheten	news,
fredrik	fredrik,
flest	most,the most,
buddy	buddy,
likaså	also,as well,
upplagan	edition,
swan	swan,
kommersiellt	commercial,
kulturell	cultural,
bli	become,
kommersiella	commercial,
köpmän	merchants,
gjordes	made,was made,
hemmet	home,
kristendom	christianity,
vasa	vasa,
åstadkomma	create,achieve,
upplysningen	the enlightenment,
kända	known,
kände	felt,
examen	exam,
disneys	disney's,
läsare	readers,
försöka	try,attempt,
chokladen	the chocolate,chocolate,
velat	wanted,
sydväst	southwest,
slogs	fought,was,
sexton	sixteen,
dagens	todays,
upp	up,
rollfigurer	roll model,role figure,
force	force,
berlins	berlin's,
förstaplatsen	first place,
bröstet	chest; breast,breast,
dennes	his,
avfall	waste,
neo	neo,
nej	no,
kommissionen	the commission,
unescos	unesco,
ned	down,bottom,
trodde	thought,
sarajevo	sarajevo,
uppdelningen	partitioning; sectionalization; division; split (-ting),division,
porträtt	portrait,
tätort	conurbation,
ort	neighborhood,place,
med	with,
genomföra	perform,
men	but,
drev	pursued,drove,led,
vinden	the wind,
mer	more,
luther	luther,
geografiskt	geographically,geographic,
därpå	darpa,thereon,
oro	worry,
åka	go,
fyllde	completed,
ajax	ajax,
sju	seven,
pilatus	pilatus,pilate,
geografiska	geographical,spatial,
dra	pull; (with)draw,
snabbast	fastest,
magnusson	magnusson,
reste	travelled,moved,
£m	million pounds,
efterföljare	following,follower,
rosenberg	rosenberg,
reagan	reagan,
atlanten	the atlantic ocean,
inleddes	started,initiated,
fördelning	distribution,
soldat	soldier,
berättelserna	the stories,tales; stories,
prokaryoter	prokaryote,
datorn	the computer,
gävle	gävle,
lennart	lennart,
provisoriska	provisional,
rockband	rock band,
oscar	oscar,
ljus	light,
nervsystemet	the nervous system,
upplevde	experienced,felt,
wikipedias	wikipedias,
ljud	sounds,
köln	cologne,köln,
kategorikvinnor	category women,
flora	flora,
trots	despite,
procent	percent,
kapitalistiska	capitalistic,
sundsvall	sundsvall,
kanadas	canada's,
erövringen	conquest,
tidskriften	the magazine,
abstrakta	abstract,
världskrigets	the world war's,
förväntade	expected,
talets	the speechs,it means "decade" but would translate as "1950s", adding an s to the year.,
klitoris	clitoris,
konstitutionen	constitution,
tusen	thousands,
tidskrifter	magazines,periodicals,
vänster	left,
satt	sat,
nobelstiftelsen	nobel foundation,
bonaparte	bonaparte,
avrättningen	execution,the execution,
trött	tired,
turnera	tour,
polis	police,
autonoma	autonomous,autonomic,
stilla	still,
orsakar	causes,
orsakas	causes,caused by,
orsakat	caused,
utomeuropeiska	non-european,
startade	started,
könsorgan	genitals,sex organ,
klarar	do,
president	president,
orsakad	caused,
indelat	divided,split,
medföra	bring,lead; result in, imply; entail,result,
indelas	divided,categorized,
indelad	divided,
medfört	resulted,
låtskrivare	song writers,
indisk	indian,
borgerliga	conservative,
kvicksilver	mercury,quicksilver,
förfäder	ancestors,
fifa	fifa,
föreställningen	the idea,the concept,
panthera	panthera,
ibrahimović	ibrahimovic,
munnen	the mouth,mouth,
murray	murray,
föreställningar	performances,notions,
helena	helena,
buddhister	budhists,buddhists,
nationell	national,
personal	personal,employed,staff,
förödande	devastating,
amerikanen	american,the american,
amerikaner	americans,
irans	iran's,
federationen	federation,the federation,
förstnämnda	first-named,aforementioned,first named,
förlängning	overtime; extension; prolongation,extension,
infektioner	infections,
aston	aston,
medlemmar	members,
downs	down,
stimulerar	stimulates,
omgivning	surroundings,surrounding,
isen	the ice,
myntades	coined,
huvudrollen	leading part,
luxemburg	luxemburg,
tillvaron	existence,the subsistence,
sida	website,side,
överraskande	surprisingly,
bröllopet	the wedding,
side	side,
kammaren	chamber,the chamber,
bond	bond,
liga	league,
päls	fur,
enorm	enormous,
medier	media,medias,
milan	milan,
aids	aids,
håret	hair,the hair,
kiev	kiev,
uppsala	uppsala,
årsåldern	age group,years old,
hänvisa	refer,
talet	rate,century,
ihop	together,
återfanns	was rediscovered,can be found,
venezuela	venezuela,
bestod	was,
foto	photo,
grundämnet	the element,element,
neutroner	neutrons,
larssons	larsson's,
normer	norms,standards,
stöds	is supported,
nietzsche	nietzsche,
nomineringar	nominations,
uppförande	construction,behavior,
folkvalda	elected,popularly elected,
faktum	fact,
iso	iso,
representant	representative,
uppbyggt	structured,
starta	startup,launch,
stewart	stewart,
gå	go,
nätet	the internet,
jordanien	jordan,
arrangeras	(is) arranged,arrange,
leddes	was led,
återkomst	return,
objektet	the object,object,
föreslagit	proposed,
girls	girls,
vikingatiden	the viking age,
förbi	past,
objekten	objects,the objects,
hollywood	hollywood,
någonstans	somewhere,
representerade	represented,
alfred	alfred,
åskådare	spectators,audience; viewer,
medeltiden	middle ages,
besegrades	defeated,
skaffade	aquired,took,
galax	galaxy,
grönwall	grönwall,
symptom	symptoms,symptom,
hundar	dogs,
formell	formal,
kontrast	contrast,
antarktis	antarctica,antarctic,
street	street,
regissören	director,
härkomst	origin,provenance,
parter	party,
troligtvis	probably,
stadsdelen	the district,district,
låta	let,
mina	my,mine,
modern	modern,
självständiga	independent,
självständigt	independent,independant,
triangel	triangle,
tecken	sign,characters,signs,
lämnar	leaves,
lämnas	left,
lämnat	left,
skildringar	scenes,description,descriptions,
tidiga	early,
monetära	monetary,
muskler	muscles,
förefaller	appear,it seems,
tidigt	at an early stage,
tål	is resistant to,stand,can take,
blue	blue,
dessa	this,these,
bildar	serves as,form,
bildas	formed; made up (of),formed,
norra	northern,
bildat	formed,
mario	mario,
luthers	luther's,
vidsträckta	wide; broad,
marie	marie,
typ	kind of,
diskuterats	been discussed,discussed,
maria	maria,
don	don,
utrustning	equipment,gear,
materiella	material,
spontant	spontaneously,
slipknot	slipknot,
vänta	(have to) wait; expect,wait,
dop	baptismal,
långvariga	long-standing,
koppla	coupling,connect,
införde	enforced,introduced,
hjälper	helps,
befälhavare	commander,
liza	liza,
droger	drugs,
skyldig	guilty,
långvarigt	long-running,long-standing,
nevada	nevada,
odling	cultivation,
krönika	chronicle,
förutsätter	assume,assumes,
folkrepubliken	people's republic,
folke	folke,
helhet	entirety,
monica	monica,
stycke	piece,piece; part; section,
meningar	sentences,
kollapsade	collapsed,
stop	stop,
stor	big; great,great,
stol	chair,
strategiska	strategical,
präster	priests,
stod	stood,
sandy	sandy,
earl	earl,
bar	bar,
bas	base,
existerar	exists,
skrivas	written,
romerskkatolska	roman catholic,
existerat	existed,
anlades	founded,were built,
fokus	focus,
förändra	change; alter; replace,change,
gärningar	deeds,
anknytning	tie,link,related,
avvikande	different,deviant; divergent; different,
zonen	the zone,
zoner	zones,
gunnar	gunnar,
vända	turn,
dittills	thus far,
vände	turned,
turnén	tour,
öppnade	opened,
inledningsvis	initially,in the beginning,by way of introduction,
skrevs	written,was,
naturligtvis	off course,naturally,
skrift	book,writing,
underart	subspecies,
göta	göta,
omkringliggande	surrounding,neighbouring,
smguld	swedish championship gold,gold medal in the swedish championships,
artikel	article,
direktör	director,
ondska	evil,
nationalister	nationalists,
harvard	harvard,
kämpa	fight,
motto	motto,
regelbundet	regularly,regularily,
isotoper	isotopes,
fns	un's,
regering	the government,
näringslivet	business,industrial life,economic life,
fördraget	the treaty,
fördragen	the compacts,
ung	young,
ernst	ernst,
regelbunden	regular,
upptäcker	discover,discoveries,
atombomberna	atomic bomb,the nuclear bombs,
gatan	street,the street,
nationalförsamlingen	national assembly,
synsättet	view,
avsikt	intention,
interna	internal,
omstritt	controversial,
varmt	warm,
erövrade	conquered,
studerat	studied,
kallats	was called,
blodkroppar	corpuscle,
cyrus	cyrus,
ting	matters,thing,
frisk	healthy,
tillämpa	administer,implement,
centralasien	central asia,
betydelsefull	meningful,significant,
igång	start,start up,
provinsen	the province,
provinser	provinces,
sällskapshundar	pet dogs,companion dog,
emigrerade	emigrated,
mindre	less,
etniskt	ethnical,
azerbajdzjan	azerbaijan,
blåvitt	blåvitt,bluewhite,blue and white,
paradiset	paradise,
ix	4,the ninth,
förgäves	in vain,
albaner	albanians,
mexico	mexico,
kvinnor	women,
ip	ip,
sushi	sushi,
dokument	files,document,documents,
in	in the context: recorded = spela (in),in,
colosseum	colosseum,
stoppa	stop,
konkurrensen	the competition,
vänstern	the left wing,left party,western,
make	husband,
producerats	produced,produced (by),
bella	bella,
västberlin	west berlin,
kommunistpartiets	communist party,the communist party,
roland	roland,
därmed	consequently,thus,
industriell	industrial,
makt	power,
benämningar	terms,names,
anglosaxiska	anglo-saxon,
atmosfären	the atmosphere,
försvarets	the defence's,
dillinger	dillinger,
skickades	sent,
kim	kim,
nicklas	niclas,nicklas,
folkrikaste	people rich,most populus,
akademiska	academical,
protesterna	protests,the protests,
roms	romes,rome's,
vetenskaplig	scientific,
sydamerika	south america,
glädje	joy,
dåvarande	then,formerly,
värmland	wermlandia,
roma	roma,
viktiga	important,
grannländer	neighboring countries,
facto	facto,
just	currently,just,
jämför	compare,
universitet	university,
psykos	phychosis,
bollen	the ball,
västeuropeiska	western european,
human	human,
anders	anders,
beskriver	describes,
premiärminister	prime minister,
fysiker	physicist,physicists,
hävdar	assert,maintain,
bokstäver	letters,
troligt	likely,
hävdat	claimed,
självstyrande	independent,self-governance,
strax	soon,just,
julen	christmas,
memoarer	memoirs,
jules	jules,
amerikas	america's,
harald	harald,
borgen	castle,the castle,
komintern	comintern,komintern,
språkets	the language's,
arkitekturen	the architecture,
gustav	gustav,
behövde	needed,
rättegång	trial,
särdrag	special features,feature,features,
följaktligen	consequently,
utrikesminister	minister of foreign affairs,
tittar	looking; viewing; viewer,
författningen	constitution,
bekräftar	confirms,
gustaf	gustaf,
trafikeras	trafficked,
trafikerar	frequent,
bekräftat	confirmed,
fastställdes	confirmed,
sjöfarten	maritime transport,
färdig	done,
medborgarskap	citizenship,
kommunerna	the municipalities,
släkting	relative,
intensiv	intense,
litauen	lithuania,
syrien	syria,
kemiska	chemical,
vattnet	water,the water,
kontinent	continent,
kunna	be able,
befolkningen	the population,
uppmärksammades	drew attention,
jupiter	jupiter,
befann	located,
kemiskt	chemically,
dominerade	dominated,
tappar	drop,lose,
statistik	statistics,
oralsex	oral sex,
miljöproblem	environmental problem,environmental problems,enviormental problem,
teoretiska	theoretical,
arthur	arthur,
däggdjuren	the mammals,
säsongerna	seasons,
shakespeare	shakespeare,
morden	murders,the murders,
filmatiserats	cinematized,screened,
mynt	coins,coin,
angrepp	attack,
burj	burj,
versioner	versions,
bolt	bolt,
härstamma	originate,
burr	burr,
förkortas	shortened,abbreviated,
super	super,
irländska	irish,
fördelen	advantage,the advantage,
ljungström	ljungström,
därutöver	in addition,moreover,
maskiner	machines,
omröstning	vote,
tolkats	interpret,interpreted,
tillverkar	makes,manufactures,
tillverkas	is made,manufacture,manufactured,
ishockey	ice hockey,
strömmar	streams,flow,
grenen	the branch,
negativa	negative,
förknippade	associated,
äktenskap	the marriage,marriage,
psykisk	psychic,
romantiska	romantic,
français	francais,public,
guide	guide,
grundades	founded,was founded,
jens	jens,
orsak	reason,cause,
utbildning	education,education and training,
havsnivån	sea level,
fastlandet	mainland,
estniska	estonian,
märks	notice,noted,
tennis	tennis,
könen	the sexes,
bönder	farmers,
bolivia	bolivia,
märke	badge,
hyllade	celebrated,
själv	alone,himself,
norrlands	northern sweden's,lapland's,
batman	batman,
sagan	story,
berg	mountain(-s),mountain,
japansk	japansk,japanese,
byggda	constructed,
bättre	better,
byggde	built,built, founded (on),
definierade	defined,
tempel	temple,
spelade	played,
positiv	positive,
slaviska	slav,slavic,slavonic,
åriga	-year,year,
regeringen	the government,government,
båten	the boat,boat,
skelett	skeleton,
månens	the moon's,the moons,
beteckningen	the label,
avsnitt	part,episode,
förändras	changes,
petit	petit,
uttryckligen	explicitly,
handelspartner	trading partner,
publiceringen	the publication,publishing,publication,
vista	vista,
handen	the hand,hand,
handel	trade,
kunnat	could have been,
svärd	sword,
betala	pay,
digital	digital,
betalt	charge,
marxism	marxism,
kungamakten	the monarchy,
överenskommelse	deal,
frodo	frodo,
exporten	the export,
accepterade	accepted,
engagemang	commitment,
riktad	directed,
ökande	increasing,
fss	fss,
expandera	expand,
riktat	pointed,
riktas	directed (at),direct,
riktar	targets,
milt	mild,
råvaror	raw,wood,raw materials,
bomben	the bomb,
telefon	telephone,
sanna	true,
manager	manager,
bomber	bombs,
vikingarna	the vikings,
marissa	marissa,
dä	with,
imperiet	the empire,empire,
avbrott	break,
uppdelning	division,partitioning,playback,
petersburg	petersburg,
dö	die,
din	yours,your,
apartheid	apartheid,
dig	up,
trenden	the trend,
afrikansk	african,
höjdes	increased,
dit	there,where,
spets	edge; top,point,
bulgarien	bulgaria,
olympia	olympia,
ville	wanted (to),wanted,
malmö	malmö,
diskografi	discography,
villa	house,villa,
slagit	beaten,
reklamen	the commercial,commercial; ad; advertisment,
invandringen	immigration,
rymden	space,
utlösning	release,ejaculation,
hästen	the horse,
bakom	behind,
afghanistan	afghanisthan,afghanistan,
viktig	important,
södra	southern,south,
föredrog	prefered,preferred,
bibliotek	library,
lennon	lennon,
somalia	somalia,
madagaskar	madagascar,
avsluta	finish,
nationalismen	nationalism,
tibet	tibet,
henry	henry,
högkvarter	head quarter,
avsaknad	absence,
kommun	municipality,
beskrivits	described,
boy	boy,
diagnoser	diagnoses,
canadian	canadian,
institute	institute,
bor	lives,
gyllene	golden,golden; gilded,
vietnamesiska	vietnamese,
mängder	amounts,
extrem	extreme,
mänsklighetens	humanity's,humanities,
hotell	hotel,
sporter	sports,
enorma	enormous,
utövar	exercise,
utövas	is practised,exercised,
världshälsoorganisationen	world health organization,
asiatiska	asiatic,asian,
sporten	the sport,sport,
religionsfrihet	freedom of religion,religious freedom,
östasien	east asia,
platån	the plateau,plateau,
franco	franco,
hemmaarena	home ground,home field,
tennisspelare	tennis player,
socialister	socialists,
semifinalen	the semi-final,semi finals,
peru	peru,
kristian	kristian,
statsmakten	the government,power,government,
österrikeungern	austria-hungary,
detaljer	details,
avsattes	dismissed,
brukade	used to,
ögon	eye (-s),eyes,
kemisk	chemical,
fartyget	vessel,ship; vessel,
fly	escape,
hände	happened,
tokyo	tokyo,
mästarna	the champions,champions,the masters,
soul	soul,
träffades	was met,reached; met,
vittnen	witnesses,
akademien	the academy,academy,riksdagens,
präglade	characterized,
anslutna	affiliated,
bristande	lack of,wanting,
sökt	searched,
ulf	ulf,
hiroshima	hiroshima,
kenneth	kenneth,
uruguay	uruguay,
winston	winston,
agent	agent,
skadades	was wounded,
utomstående	outside people; outsiders,outsider,
dennis	dennis,
kunglig	royal,
pink	pink,
diskuterades	discussed,
oslo	oslo,
engelsmännen	english people,the english,the british,
återvänder	returns,
ekonomiska	economical,
till	to,
gitarrist	guitarist,
nya	new,
nye	new,
mat	food,
regeringstid	term of government,term of government; term of office,reign,
may	may,
överensstämmer	conform,agree,match,
uppföljare	sequel,
fotboll	football,
läkare	doctors,doctor,
maj	may,
upphört	ceased,
man	one,
asien	asia,
johnson	johnson,
sådana	such,
q	q,
tala	speak,
block	block,
basket	basketball,
romantiken	romance,romanticism,
undantag	exception,
sådant	such,
lsd	lsd,
bussar	bus,
bevisa	prove,
alfabetet	the alphabet,
unionen	union,the union,european union,
gällde	applied,applied to,
sällsynta	rare,
moralisk	moralic,moral,
huvudsak	in principal; chiefly,mainly,main thing,
lyrik	poetry,
motståndet	the resistance,the resistence,
verksam	active,effective,
landskap	province,landscapes,landscape,
juryn	the selection panel,the jury,
sekter	sects,
inkomster	income,
äkta	genuine,married,authentic,
nazisterna	the nazis,nazis,
policy	policy,
växte	grew,grow,
main	main,
texas	texas,
lägst	lowest,lowermost,
steget	step,
janeiro	janeiro,
domstolar	courts,
försörjning	sustention,sustentation,
sibirien	siberia,
leds	led by,passed,
vindkraft	wind power,wind,
färg	colors,colour,
uppskattning	appreciation,estimated,
leda	lead,
villkoren	the terms,conditions,
fortsättning	continuation,
tysklands	germany's,germanys,
latin	latin,
tacitus	tacitus,
sökte	searched,
söner	sons,
vattendrag	streams,watercourse,
avkomma	offspring,
dianno	di'anno,dianno,
saudiarabien	saudi arabia,
canada	canada,
jackson	mrs. jackson,jackson,
håkansson	hakansson,
avrättningar	execution,executions,
pamela	pamela,
områdena	the areas,areas,
tronföljare	heir,successor,
kattdjur	felidae,cat,
valdes	chosen; elected,
premiären	premiere,premier,
monster	monster,
romani	romany,roma,
konstnär	artist,
chiles	chile's,
tomt	empty,
dubbla	double,
california	california,
miley	miley,
brooke	brooke,
kognitiva	cognitive,
ord	word,words,
tunnelbanan	subway; tube; underground,the subway,
keith	keith,
verkade	did,were active, worked, was active,
gott	practically; good,
anledning	reason,
självmord	suicide,
uppvisar	shows,
rankningar	ranking,rankings,
vision	vision,
stängdes	closed,
kraftig	strong,
egentligen	actually,
centrala	central,
grupperna	groups,
intryck	impression,
uttalanden	statements,
här	this; here,is,here,
rachel	rachel,
folklig	popular,
centralt	central,
skapandet	creation,the making,
kommunism	communism,
sätt	manner,way,
homogen	homogenous,
visar	shows,
består	consists of,exists,
västbanken	the west bank,westbank,
grundämnen	elements,
individ	individual,
örebro	Örebro,
öronen	the ears,
besluten	decisions,
anus	ass,anus,
köpenhamns	copenhagen's,
fysiska	physical,
fysiskt	physically,physical,
danny	danny,
löstes	solved,
drevs	concentrated,was driven,
beslutet	the decision,
konkreta	concrete,
fiender	enemies,
fienden	the enemy,
medlemmarna	the members,
lugn	calm,
sean	seab,
fordon	vehicle/-s,vehicles,vehicle,
inträde	entry,
marklund	marklund,
jämlikhet	equality,
stadsdelar	districts,city districts,
större	bigger,
formerna	forms,
tänder	teeth,
orsakerna	the causes,
kevin	kevin,
adeln	nobility,
nikola	nikola,
politiska	politic,
förälskad	in love,
menas	means,
skulptur	sculpture,
centralbanken	centralbank,central bank,
potential	potential,
politiskt	political,
performance	uppträdande,
centralstation	central station,
magnetiska	magnetic,
channel	channel,
norman	norman,
isolerad	isolated,
hertig	duke,
livets	life's,the life's,
halvan	the half,half,
politisk	political,
teoretiskt	theoretic,theoretical,
mordet	the murder,
beskrivit	described,
civilisationer	civilizations,
visades	showed,
otaliga	countless; endless,countless,
lojalitet	loyality,loyalty,
drottning	queen,
grammatik	grammar,
österut	eastwards,east,
kontrolleras	is controlled,
kontrollerar	controlling,controls; controlling,
ungdom	youth,
civilisationen	civilization,
adolfs	adolf's,
uranus	uranus,
tidigast	the earliest,
samlingsalbum	compilation album,
helig	holy,
dick	dick,
historier	stories,history,
passande	fitting,suitable,
historien	history,
black	black,
medeltidens	medieval,
lyssnade	listened,
ges	given,be given,
ger	gives; is giving,give,
raser	species,
kulturellt	cultural,culturally,
motsvarande	corresponding,
ramadan	ramadan,
landets	the country's,
katla	katla,katla (fictive dragon in the classic "bröderna lejonhjärta"),
vintergatan	milky way,the milky way,
firade	celebrated,
ledaren	leader,
gen	gene,
rasen	the race,
himmlers	himmlers,
mattis	mattis,
bengtsson	bengtsson,
statistiska	statistical,
förenta	united,
spridda	spread,scattered,
världskrigen	the world wars,
europacupen	euro (-pean) cup,european cup,
london	london,
tolfte	twelth,
relativt	relatively,
sämre	poor,
hittar	finds,
fokuserar	focuses,focus,
toppade	topped,
relativa	relative,
jordytan	earth crust,
slöt	joined (in peace),closed,
utgiven	published,
menat	meant,
menar	means,
kandidater	candidates,
försvarsmakten	national defense,national defence,
döden	death,
vanns	(was) won,
människan	the human,
söndagen	sunday,
personligt	personal,
världskriget	world war,
gaga	gaga,
människas	human's; man's,human,
personliga	personal,
tsaren	the czar,the tsar,
august	august,
ju	the,the more,
tur	turn,
forskaren	researcher,
jr	junior,
åker	go,field; going,
timme	hour,
tum	inch,
signaler	signals,
lexikon	lexicon,
ja	yes,
ministrar	ministers,
rugby	american fotboll,rugby,
ån	on,the river,
utvalda	selected,selected; chosen,
tour	tour,
åt	to,for,
ås	ridge,site,
år	the year,
vätska	fluid,liquid,
naturresurser	natural resources,
tryck	print,pressure,
väst	west,the west,
århundraden	centuries,
cancer	cancer,
statschefen	the head of state,
syntes	synthesis,
mariette	mariette,
grundare	founder,
territorium	territory,
mätningar	measurements,
ryggen	the back,
barry	barry,
överföra	transfer,
bildats	had formed,created,
kirsten	kirsten,
industrin	industry,
västliga	western,
mars	march,
överförs	transfered,
plötsligt	suddenly,sudden,
marx	marx,
mary	mary,
kultur	culture,
handels	trade,
flaggan	the flag,
cobain	cobain,
partido	partido,
avskaffa	abolish,
bmi	bmi,
jagar	hunts,hunting,
spelfilmer	motion pictures,feature film,feature films,
skrivet	written,
fortsatt	continued,
metall	metal,
dragit	drawn,dragged,
uppstod	developed,
kategorimän	category: men,
insåg	realized,
nionde	ninth,
sahara	sahara,
däribland	among them,including,
uppmanade	urged,encouraged,
liknande	similiar,similar,
uppfyller	fulfills,
hålls	is held,maintaned,
par	pair,
upplagor	the edition,issues,
jesu	jesus,
beredd	ready (to),prepared,
lava	lava,
hålla	keep,
röka	smoke,
stött	met,
samt	also,as well as,
hösten	the fall,the autumn,
kuba	cuba,
teknisk	technical,
lösningar	solutions,
sömn	sleep,
markus	marcus,
gates	gates,
münchen	munich,
bebyggelse	settlement,settlements,habitation,
reaktionen	the reaction,
dinosaurierna	dinosaurs,
byggnad	building,
reaktioner	reactions,
våld	violence,
jakten	the hunt,
ideologiskt	ideological,
grannländerna	neighbouring countries,
avskaffandet	abolition,abolishment,
programledare	host,
gotland	gotland,
ideologiska	ideological,
motverka	prevent,counteract,counter,
trä	wood,
hanen	the male,
vintern	the winter,winter,
schwarzenegger	schwarzenegger,
underarten	subspecies,sub species,
mån	mon,
mor	mother,
haft	had,
prägel	mark,
mot	against,
kategori	category,
jakt	hunt,hunting,
simmons	simmons,
underarter	sub-species,subspecies,
baltiska	baltic,
kollektiv	collective,
mod	courage,
christina	christina,
adams	adams,
började	started,began,
födde	gave birth too,
jordbävningar	earthquakes,
manhattan	manhattan,
mänsklig	human,
sågs	seen,was observed,
göran	göran,
bipolära	bipolar,
göras	made,be made,
grannar	neighbours,
joan	joan,
feodala	feudal,
maos	maos,mao's,
förs	led,
jordbruket	the agriculture,
lotta	lotta,
fört	led,lead,
sudan	the sudan,
reportrar	reporters,
föra	pre,lead,
före	ahead (of), before,before,
ända	as far as,
demokratisk	democratic,
traditionell	traditional,
ände	end,
moderata	moderate,moderates,
vistas	live,present,
förlust	loss,
londons	london's,
cellen	the cell,
olof	olof,
akon	akon,
tongivande	influential,
tillverka	producing,
sjätte	sixth,
celler	cells,
allians	alliance,
metaforer	metaphores,metaphors,metafor,
lands	on land,
lagarna	the laws,
retoriken	rhetoric,
herbert	herbert,
newtons	newton's,
wilde	wilde,
dödsfall	death,
mark	ground, soil, territory,ground,
intellektuella	intellectuals,
floderna	floods,the rivers,
fullständigt	completely,
gravid	pregnant,
behandling	treatment,
varelse	creature,
emellanåt	once in a while,occasionally,
anfalla	attack,
välmående	well-being; affluent,prosperous,
fullständiga	complete,
kvinnlig	female,
tillfälligt	temporarly,temporary,
eget	own,
inletts	started,
utbredd	widespread,
birger	birger,
härifrån	from here,
e	e,
egen	own,
tävlingen	competition,contest,
vhs	vhs,
exemplar	copies,
bibliografi	bibliography,
manuel	manuel,
verkliga	real,
kröntes	been crowned,crowned,
humanismen	humanism,
parlament	parliament,
följde	followed,
youtube	youtube,
manliga	male,
öns	the islands,island's,
prestigefyllda	prestigious,
skriven	written,
pompejus	pompey,pompejus,
arabiska	arabic,arabian,
goebbels	geobbels,
film	film,
genrer	genres,
effekt	effect,
istanbul	istanbul,
spåren	the tracks,tracks,wake,
rubiks	rubik's,
muren	wall,
produktiv	productive,
stannade	stayed,
faktorer	factors,
däremot	on the contrary,however, on the contrary,
ordna	arranging,arrange,
profet	prophet,
ungarna	the kids,the young,
ledning	guidance,
kyros	cyrus,
världsliga	worldly,
medicinska	medicinal,medical,
araberna	arabs,
palestinska	palestinian,
uppfostran	upbringing,
medicinskt	medical,
god	good,
snabbaste	fastest,
begå	commit,
resolution	resolution,
åtskilda	segregated,separate,
vila	rest,
socialismen	the socialism,socialism,
inspirerat	inspired,
dollar	dollar,
vill	will,want,
hindrar	prevents,stop; prevent,
ingripande	intervention,
inspirerad	inspired,
levern	the liver,
zink	zinc,
symbolen	the symbol,
lugna	reassure,calm,
rwanda	rwanda,
symboler	symbols,
skydda	protect,
skriver	write,
seriens	series,
kasta	throw,
avhandling	thesis,
handlade	dealt with,was (about); traded,
israeliska	israeli,isrealic,
ramen	frame,
stödja	support,
ramel	ramel,
kulminerade	culminated,
ansvarig	charge,
miljoner	millions,
båtar	boats,
snuset	snuff,the snuff,
suttit	sat,
massor	lots,(in) masses,
växthuseffekten	the greenhouse effect,greenhouse effect,
intressant	interestingly,
material	material,
abc	abc (swedish news program),
danmark	denmark,
publik	audience,public,
östtysklands	east germany's,
lärare	teacher,
värderingar	evaluations,
långhårig	long-haired,
bebott	inhabit,inhabited,an inhabitated,
närhet	proximity,closeness,
vald	elected,
jonas	jonas,
benen	legs,
valt	chosen,
sångare	singer,
historiker	historians,
uppslagsverk	encyklopedia,
alexandria	alexandria,
sjukhuset	the hospital,
africa	africa,
enat	united,
rösterna	votes,the votes,
författaren	the author,
hyllning	tribute; homage,
torrt	dry,
utmärkelsen	award,the award,
innebar	meant,was; meant; entailed,
utmärkelser	commendations,awards,
torra	dry,
landet	state,the country,
diamond	diamond,
människa	man,
romersk	roman,
koma	coma,
brist	lack,failure; lack of,
tillkommer	reside,will be added,
hundraser	breed of dogs,
skivor	records,
berätta	tell,
flytt	escaped,fled,
tillverkningen	production,the production,
det	it,
roosevelt	roosevelt,
utsläpp	emissions,
bron	the bridge,
del	part,
lindgren	lindgren,
lagerlöf	lagerlöf,
baháulláh	bahullah,
befintliga	existing,
samtliga	all,
hastigt	fast,
latinets	the latin,the latin's,
sovjetunionens	soviet union's; soviet's,
hjälpte	helped,
sjukdom	illness,disease,
medförde	resulted,brought,led,
födseln	the birth,
sträng	string,
robinson	robinson,
protein	protein,
makten	the power,
hämta	fetch,
psykotiska	psychotic,
georgien	georgia,
stig	stig,
verkligheten	reality,
blad	leaves,leaf,
försvinner	disappears,disappearing,disappear,
primära	primary,
vikten	importance,
makter	powers,
rastafari	rastafari,rastafarian,
avtalet	the treaty,the contract,
pettersson	pettersson,
laboratorium	laboratory,
huvudkontor	central office,headquarters,
ligger	lies,is,
vatten	water,
rastafarianer	the rastafarian,rastafarian,rastafarians,
rockgrupper	rock groups,rock group,rock bands,
facebook	facebook,
paz	paz,
konservatismen	conservatism,
civila	civil,
inåt	inwards,
nordsjön	north sea,
officiella	official,
latinamerika	latin america,
fältet	the field,field,
höll	held,hold,gave,
göra	do,do; doing,
försäkra	insure,make sure,assure,
tvåa	second,
same	lapp,
görs	made,is made to,
officiellt	officially,
människans	humans,mankinds,
längden	lenght,
diskussion	discussion,
wilhelm	wilhelm,
edmund	edmund,
inbördeskriget	civil war; civil war,civil war,
epok	epoch,
gustafsson	gustafsson,
saknades	lacked,missing,
trossamfund	religious community,faith community,
suverän	terrific,supreme,
träffar	meets,
ställas	set,be set,
planerna	the plans,
fängelse	prison,
sexuellt	sexual,
oxford	oxford,
skrifterna	scriptures,
porto	postage,
robbie	robbie,
kungarna	the kings,
namibia	namibia,
inleder	initiates,
haile	haile,
mental	mental,
fisk	fish,
flytta	move,
öron	ears,
förenade	united,
energi	energy,
perry	perry,
sanningen	the truth,
östman	Östman,
oftast	usually,most often,
infrastrukturen	infrastructure,the infrastructure,
ölet	the beer,
forskning	research,
perro	perro,
förföljelser	persecution,pursuits,persecutions,
fullständig	n/a,
konflikt	conflict; strife,
bränslen	fuel,
lawrence	lawrence,
strömning	flow,
eventuella	eventual,
blekinge	blekinge,
uralbergen	the ural mountains,
eventuellt	eventually,possibly,
helsingör	helsingör,
inflationen	inflation,
legender	legends,
finland	finland,
styrs	ruled,
fått	was given,
styre	rule,
legenden	legend,
ensam	alone,
styra	steer,
top	top,
sjunkande	sinking; decreasing,
säkerhetsråd	security council,
treenighetsläran	doctrine of the holy trinity,trinity,school of trinity,
snarast	rather,as soon as possible,
juridiska	juridical,legal,
carter	carter,
kom	came,
kol	coal; charcoal,
gator	streets,
åtta	eight,
observationer	observations,
förhindrar	prevents,
kardinal	cardinal,
järnvägar	failways,railways,
triangeln	the triangle,
gudarna	the gods,
domstolen	the court,
början	beginning,
matteusevangeliet	gospel of matthew,book of matthew,
följden	the result,the cause,result,
fort	quickly,
b	b,
knapp	scarce,bare,
proteinerna	the proteins,
ö	island,
personens	the persons,the person's,
singapores	singapores,singapore's,
hellström	hellström,
baháí	bahá'í,
avtar	declines,
självständig	independent,independant,
följder	consequences,
följdes	followed,was followed,
rikedom	riches,wealth,
försökte	tried to,tried,
bränsle	fuel,
gjord	made,
adjektiv	adjective,
gjort	made,created,
hundratals	hundreds of,hundreds,
stewie	stewie,
mussolini	mussolini,mossolini,
infrastruktur	infrastructure,
caesar	caesar,
genast	at once,
taktik	tactics,tactic,strategy,
inkomsterna	the incomes,
dramatiskt	dramatically,
skjuta	postpone; shoot,
varifrån	from where; wherefrom,from which,
patterson	patterson,
krafter	forces,
gillade	liked,approved; liked,
niclas	niclas,
kraften	the force,
utbrott	outbreak,
samtidigt	simultaneous,
laila	laila,
högt	high,
ko	cow,
km	kilometers,
kl	hr,o'clock,
höga	high,
organisk	organic,
organism	organism,
thomas	thomas,
venedig	venice,venedig,
kvalitet	quality,
gradvis	gradually,
relation	relation,
utveckla	develop,developing,
fina	fine,
nämns	mentioned,
antagit	presumed,
konto	account,
undre	lower,
wallenberg	wallenberg,
medverka	take part,participate,
världens	the world's,the worlds,
tionde	tenth,
religionerna	religions,the religions,
förbudet	the union,
avseende	regard,
blomstrade	flourished,
typiskt	typical,
notation	notation,
beslutar	decides,
vänskap	friendship,
express	express,
beslutat	resolved,decided,
förklarat	explained,declare,
typiska	typical,
husen	the houses,
skickas	is sent,sent,
skickar	sends,send,
brukar	usually,used to,
wallander	wallander,
bindande	binding,
uttrycket	the expression,
uttrycker	express,express (-es),
huset	the house,
somrar	summers,
stadium	stage,
styrdes	was guided,governed,ruled,
suveränitet	sovereignty,
rollfigur	character,
godkännas	pass on,be approved,
höglandet	highlands,the highland,
händelsen	the occurence,event,
fann	found,
rovdjur	predator,
fans	fans,
landsbygden	rural area,
champagne	champagne,
romarriket	the roman empire,
bildandet	setting-up,establishment,
professionella	professional,
framförs	is presented,
framfört	expressed,presented,
rörelserna	the movements,
kritiserades	critisized,
framföra	convey,
skivorna	the records,records,
medlem	member,
musklerna	the muscles,
statligt	state,governmental,
vuxit	grown,
restaurang	restaurang,
baltimore	baltimore,
romska	romani,
beta	graze,
globala	global,
kroatiens	croatia's,croatias,
förklaring	explaination,explanation,
point	point,
folkmord	genocide,
karaktären	the character,character,
andas	breath,
orsaken	reason,cause,
således	hence,thus,
tennessee	tennessee,
globalt	globally,
behöll	kept,
våningar	floors,storeys,
laos	laos,
fördrevs	was banished,driven away,
konspirationsteorier	conspiracy theories,
inför	before,
bengt	bengt,
popularitet	popularity,
gav	gave,
effektiva	effective,
gas	gas,
vana	familiar,used,habit,
kalmar	kalmar,
effektivt	effective,
trupperna	the troops,
detsamma	the same,
bild	picture,
motorväg	freeway,highway,
åtalades	was prosecuted,charged,
spridning	diffusion,distribution,
döptes	renamed; named,renamed,baptised,
portugal	portugal,
arenan	arena,
elektronik	electronics,
påbörjade	started,
monroe	monroe - it's a persons name,monroe,
rederiet	the shipping company,the company,shipping company,
dödat	killed,
granska	review,
sjuk	ill,
dödar	kills,
dödas	put to death,killed,
hamna	end up,
tänkt	supposed; intended,intended,
administrationen	administration,
tyder	indicates,
sapiens	sapiens,
övertogs	overtaken,
skotska	scottish,
syd	south,
syn	view,
jerusalems	jerusalem's,
koloniala	colonial,
avsett	regard,intended,
nämnde	mentioned,
småningom	when the time comes,eventually,
tillbehör	sides,condiments,accessory,
nämnda	said,
kungariket	kingdom,the kingdom,
noll	zero,
kapitel	chapter,
albanien	albania,
regim	regime,
ministerrådet	minister counsellor,
värme	heat,
skott	bulkheads,round,shots,
halva	half,
norrland	norrland,
dikter	poems,
bibeln	bible,
kommunister	communists,
juventus	juventus,
halvt	half,
verkställande	executive,
passerar	passes,
struktur	structure,
senaste	last,
alternativt	alternatively,alternative,
analytiska	analytical,
alternativa	alternative,
tropisk	tropical,
sektion	section,
sparta	sparta,
administrativt	administrative,administratively,
monarkin	the monarchy,
dömd	sentenced,convicted,
administrativa	administrative,administative,
åtal	prosecution,
dubbelt	double,
bil	car,
teknik	technique,technology,technic,
big	big,
kejsaren	the emperor,
avlidna	the perished,
möttes	met,
bit	piece,
indonesiska	indonesian,
situationen	situation,the situation,
rené	rené,
grå	gray,grey,
kolonialtiden	the colonial times,
princip	principle,principal,
möjlig	possible,
stränga	severe,
tillstånd	to the dental,condition,
anatomi	anatomy,
google	google,
identisk	identical,
egyptiska	egyptian,
tolkningar	interpretations,interpretation,
verkat	worked,acted,
studerar	study,studies,
cocacola	coca cola,coca-cola,
lars	lars,
västergötland	västergötland,
flygplatser	airports,air ports,
måste	have to,
integration	integration,
per	per,
pratar	talking,talk,
självstyre	self-governance,
energin	the energy,
lösningen	the solution,solution,
därför	because,therefore,
nordamerika	north america,
resande	travelling,
påven	the pope,
ockuperade	occupied,
britannica	britannica,
korta	short,
värmestrålningen	heat radiation,
uppfattningar	opinions,
fallit	fallen,
jimmy	jimmy,
grammy	grammy,
styrelse	government; direction,board of directors,
barcelonas	barcelona's,
steven	steven,
ordnar	fix,decorations,arrange,
brita	brita,
ontario	ontario,
framträdde	appeared,
ökningen	the increase,
ansvar	responsibility,
turkiska	turkish,
medvetande	consciousness,awareness,
jaga	hunt,chase,
serie	comic; row; succession; serial,cartoon,
konsul	consul,
bostäder	residences,
torsten	torsten,
jonathan	jonathan,
skillnaden	the difference,
lånat	borrowed,
mångfald	diversity,variety,
planet	planet,
smycken	jewlery,
sultanen	sultan,
planer	plans,
reggaen	the reggae,
jordbävningen	the earthquake,
reidar	reidar,
titel	title,
expedition	expidition,expedition,
förbjudna	forbidden,prohibited,
hjärnans	the brain's,
tropiskt	tropical,
tropiska	tropical,tropic,
materia	materia,
tyskland	germany,
eller	or,
voltaire	voltaire,
familjer	families,
årstiderna	the seasons,
familjen	the family,
betalar	pay,
makedonien	macedonia,
anser	believes,
anses	deemed; regarded,
förr	sooner; past,sooner,
lena	lena,
utvecklade	developed,
länders	countries',countrie's,
samla	gather,
mutationer	mutations,
nådde	reached,
ritualer	rituals,
talades	spoken,spoken (of),spoke,
sambandet	the connection,connection,relation,
dramatiker	dramatists,
förbjudet	prohibited,
judisk	jewish,
öppnat	opened,
regionalt	regional,regionally,
flod	river,
stänga	close,
stred	fought,
frankrike	france,
förut	before,
sigmund	sigmund,
stängt	closed,
intensivt	intensive,
privat	private,
tillämpningar	situations,implementations,
medlemskap	membership,
betrakta	view; regard,view,
sydafrikanska	south african,
sahlin	sahlin,
konsten	art,the art,
intensiva	intensive,intense,
kollaps	collapse,
atlas	atlas,
protokoll	protocol,
nobelpriset	the nobel prize,
luleå	luleå,
kampanjen	campaign,
turkiets	turkey's,turkeys,
annika	annika,
tjänade	earned,
varnade	warned,
utgjordes	make up,comprised; consisted,
tävlingar	competitions,contests,
exemplet	the example,example,
knight	knight,
joel	joel,
samman	together,
slutade	quit,
vanligen	usually,
warszawa	warzaw,warsaw,
endast	only,merely,
joey	joey,
tunnlar	tunnels,
störtades	overthrew,overthrown,was overthrown,
överhöghet	supremacy,suzeranity,sovereignty,
utbredda	widespread,
vanligaste	frequent,most common,
påsken	easter,
earth	earth,
depression	depression,
sträcker	stretches,
går	goes,
chicago	chicago,
tillkomst	established,
effekter	effects; repercussions,
sauron	sauron,
placering	placement,
vätet	the hydrogen,
och	and,
kyrka	church,
öar	islands,
extremt	extreme,
ordförande	chairman,
börja	start,
extrema	extreme,
isländska	icelandic,
befolkningstäthet	population density,
populäraste	most popular,
sina	their,
honom	him,
svårigheter	difficulties,hardships,
medeltid	the medieval times,
skada	damage,
alaska	alaska,
katolicismen	catholisism,
lagförslag	bill,
miljard	billion,
honor	ära,
färgade	colored,
existens	existence,
uppnår	achieve,
uppnås	is achieved,
talare	speaker,spoke,
privata	private,
stundom	sometimes,somtimes,
når	reach,
nås	reached,
filippinerna	the philippines,
betraktar	regard,
nåd	mercy,
lima	lima,
somrarna	the summers,
skivbolag	record company,
kinesisk	chinese,
skotsk	scottish,
chi	chi,
gruppspelet	groupplay,group play,
fånga	capture,
döpt	named,baptized,
linköpings	linköping's,
nytta	good,useful,
geografisk	geographic,geographical,
titanics	titanic's,
iis	ii's,
prinsen	prince,the prince,
platser	places,
utropade	cried out,
bakterier	bacteria,
självständighet	independence,
avsikten	intention,
iii	iii,
platsen	the place,
ansvaret	responsibility,the responsiblity,
britney	britney,
f	f,
tunnel	tunnel,
påbörjas	starts,begin,
arton	18,eighteen,
baserad	based,
kedja	chain,
kategorisvenska	category: swedish,
baseras	based,bases,based on,
baserar	based,
baserat	based,
kyrkan	the church,
väldet	empire,the rule,
fotosyntesen	photosynthesis,
titlar	titles,
mozarts	mozart's,
cecilia	cecilia,
fett	fat,
internationellt	international,internationally,
lanserade	introduced,
internationella	international,
vilhelm	vilhelm,
revs	was demolished,
böckerna	books,
rousseau	rousseau,
riktig	real,
klar	done,
expansionen	the expansion,
malta	malta,
föddes	was born,born,
herrlandskamper	men's international contest,men's international contests,
brändes	burned,
spannmål	grain,
förbundskapten	manager,coach,
klan	clan,
gammal	old,
terrier	terrier,
siv	siv,
finländska	finish,finnish,
rådhus	courthouse,
dryck	drink,drinks,
förekommit	occured,
billboardlistan	bilboardlist,
registrerade	noted,
olyckan	the accident,
alltjämt	remains,
bilbo	bilbo,
omslaget	the cover,
meter	metre,meter,
strid	fight,
innebär	mean,means,
le	smile,
människor	people,
la	la,
variationer	variations,
bryts	breaks,
tvungna	forced,forced to,
tillägg	addition,
weber	weber,
dag	dag,day,
spektrum	spectra,spectrum,
utfärdade	issued,
slags	kind,
dam	dam,lady,
valet	the election,
tillkommit	accured,
periodiska	periodic,
sammanhanget	context,
installera	installing,install,
day	day,
kontinuerligt	continuous,continous,
beslut	decision,
februari	february,februari,
syftade	alluded to,aimed,
lysande	brilliant,
engelskspråkiga	the english language,
juridisk	legal,
krita	chalk,
humanism	humanistic,humanism,
kristiansson	kristiansen,
dokumentär	documentary,
inspirerade	inspired,
segern	the victory,
marley	marley,bob marley = singer,
arbetskraft	labor,
fattigdomen	poverty,
nödvändiga	essential,
matt	matt,
jerusalem	jerusalem,
mats	mat's,
kärnan	core,
nödvändigt	necessary,
deras	their,
upphörde	ceased,expired,discontinued,
återta	retake,regain,reclaim,
webbplats	website,
franz	franz,
odlas	cultured,
arbetare	workers,
längre	longer,
inleds	starts,
efterträddes	succeeded,
medelhavsområdet	the mediterranean region,the mediterranean area,
farbror	uncle,
fotografier	photographs,
nivå	level,
south	south,
liberaler	liberals,
stämmer	(if it's) true,is true,
genomgår	undergoes,undergoing,
pga	because of (short of "på grund av"),
uppger	states,
innehålla	include,contain,
insikt	insight,recognition,
levnadsstandarden	the standard of living,living standard,
fruktade	feared,
omständigheter	circumstances,
veckan	the week,
leder	leads,leading (to),
utlopp	outflow,
energikällor	energy resources,energy sources,sources of energy,
kantonerna	the cantons,cantons,
förklara	explain,
leden	lines,the route,
palestina	palestine,
demonstrationer	demonstrations,
bundna	bound,tied,
noterade	noted,
stället	instead,the place,
ställer	running; causing,run (in election),
innehade	possessed,
firades	was,was celebrated,
utföra	perform,
ledamöter	commissioners,
släkten	the family,
ställen	spots; places,places,
bevarats	protected,preserved,
beskrivningen	description,
domaren	the judge,
matematisk	mathematical,mathematic,
uteslutande	exclusivly,
osmanska	osmanian,ottoman; osmanli,
universum	universe,
mälaren	mälaren,
premiär	premiere,
havs	at sea,
aristoteles	aristoteles,
biologiska	biological,
operativsystem	operating system,
följd	effect,
älgar	moose,
följa	follow,
basist	bassist,
uganda	uganda,
idag	today,
rådande	current,prevalent,
följt	followed,
mil	mile,swedish miles,
min	my,
fötter	feet,on its feet,
kroppar	bodies,
tidningar	magazines,
mig	me,
låg	low,
experter	experts,
lån	loan,
konstverk	work of art,artwork,
konkurrerande	competing,
framförts	performed,
resurser	resources,
resultatet	the result,result,
dinosaurier	dinosaurs,
varandras	each others,each other's,
missionärer	missioners,missioner,
resultaten	the results,
sedan	since,
sist	last,
herman	herman,
liknade	looked like,
stranden	shore,the beach,
republikanska	republican,
rörelsens	operating,movements,
milano	milano,
deuterium	deuterium,
tidskrift	newspaper,magazine,
capita	capita,
styrke	strength,been,
definiera	define,
viktigaste	most important,
styrka	strength,
utgångspunkt	starting point,point of departure,
högtider	holiday,
text	text,
charles	charles,
inhemsk	domestic,native,
ugglas	ugglas,
timmar	hours,
kurfursten	elector,
rumänska	romanian,
järnvägen	railroad,
euroområdet	eurozone,
rytmiska	rhythmic,more rhythmic,
temperatur	temperature,
satan	satan,
shahen	the shah,
säker	safe,
bryssel	brussels,
organiska	organic,
snitt	on average,average,
influensavirus	flu virus,flue virus,
förändrades	changed,
buddhismen	buddism,buddhismen,
överlägset	superior,
förstår	understand,
regimen	regime,
studenterna	the students,
uppehåll	pause,hiatus,
vinsten	the win,
organ	body,agency,organ,
nazitysklands	nazi germany's,nazi germany,
vinster	profit,
majoriteten	the majority,
lyckade	successful,
byggdes	was built,
ronaldo	ronaldo,
svenske	swedish,
svenska	swedish,
eleonora	eleonora,
kapitalet	the capital,
först	first,
egentlig	actual; factual; real,actual,
reform	reform,
redan	already,has already,
konverterade	converted,
ordnade	arranged,
bruno	bruno,
avslutades	ended; concluded,concludes,
bör	should,
ordentligt	proper,properly,
översikt	overview,
koncept	concept,
industrialisering	industrialization,
uppskattade	appreciated,
listan	the list,
hårdare	harder,more severely,
säkerheten	the security,
översättas	translated,translated (to),
viktigare	more important,
läsning	reading,
hämtade	brought,
buddhas	buddha's,
konservativa	conservative,
miniatyr|karta	miniature|map,
återförening	reunion,
litteratur	litterature,
aktuellt	current,
förekommande	occuring,
kommunicerar	communicates,
regimer	regimes,
aktuella	current,
kommendör	commandor,commander,
sachsen	saxony,
fester	parties,
inneburit	meant,
befogenhet	warrant,authorization,authority,
utsågs	appointed,was appointed,
medicinsk	medical,
elektroner	electrons,
ad	ad,
af	of (old swedish),
grupperingar	groups,groupings,
slippa	avoid,
gaza	gaza,
igen	again,recognize,
asteroider	astroids,asteroids,
försvar	defence,
stationen	station,
stationer	stations,
orange	orange,
västmakterna	western powers,
uppmärksammat	noticed,
general	general,
napoleon	napoleon,
augusti	august,
bruket	the use,
kraftiga	powerful,
stalin	stalin,
ar	is,
ocheller	and/or,
betraktade	considered,
palats	palaces,
tagits	taken,
flyktingar	refugees,
verkligen	real,the reality,
fördrag	agreement,treaty,
vistelse	visit,stay,
prosa	prose,
utom	except,
händelserna	the events,the happenings,
lämnade	left,
wolfgang	wolfgang,
blodtrycket	blood pressure,
sångerna	song are,the songs,
omedelbart	immediately,
heinrich	heinrich,
hinduismen	hinduism,up,
kallad	called,
kontrollera	control,
framförallt	above all,in particular; above all,
kallat	called,
kallas	called,
kallar	calls,
center	center,
thailand	thailand,
seth	seth,
antonio	antonio,
sett	seen,except,
hoppas	hope,
omgångar	in turns; periods; mandates,
svensk	swedish,
undvika	avoid,
deltar	participates,
stores	the great's,the great,
kontaktade	contacted,
passade	suiting,fit; suited,
mystiska	mystical,
wagner	wagner,
misshandel	abuse,
grekiskans	the greek's,greek,
flertal	several,majority group,
vanligt	usual,
hamburg	hamburg,
kampf	on,kampf,
liverpools	liverpool's,liverpools,
reformer	reformers,reforms,
anhöriga	relatives,
lake	lake,
mentala	mental,mentala,
landområden	land,land areas,
streck	bar,
match	game,match,
förnuft	common sense,reason,
uppmärksamhet	attention,attantion,
uppträder	appears,performs,occur,
dubai	dubai,
demens	dementia,
innehöll	include,
chrusjtjov	chrusjtjov,
viruset	virus,
likt	like,
journalist	journalist,
uppträda	appear,act,
gudomlig	divine,
albumets	album's,
starkaste	strongest,the strongest,
insats	contribution,intermediate,stake,
etablerades	was established,
minsta	minimum,
joachim	joachim,
löser	solves,
skildrar	describes,
skildras	is depicted,depicted,
gisslan	hostage,
internationalen	international,
definitionen	definition,the definition,
nattetid	overnight,
definitioner	definitions,
starkare	stronger,
leopold	leopold,
arterna	the species,
nordkorea	north korea,
socker	sugar,
ärkebiskopen	archbishop,
glada	happy,
mäktigaste	powerful,most powerful,
slutgiltiga	final,
andel	share,
anden	the holy spirit,
folkräkningen	census,
medverkar	contribute,
alexanders	alexanders,alexander's,
rörde	was about,
socken	parish,
omgiven	surrounded,
potatis	potato,
tränger	forces forward,cut in,
skapade	made,created,
australiska	australian,
ljusare	brighter,lighter,
föredrar	prefer,
vimmerby	vimmerby,
hatar	hate,hates,
densamma	the same,
skog	forest,
kuben	the cube,
strävhårig	hispid,wirehaired,
föga	little,hardly; little,
kärnor	cores,
kväll	evening,
klockan	clock,o'clock,
civilbefolkningen	civilian population,the civilian population,
ryssarna	the russians,
brand	fire,
bröder	brothers,
ersättning	pay,
flygvapnet	air force,the airforce,
kraft	force,power,
bud	bid,message,
vetenskap	science,
utrymme	space,
arbetsgivaren	employer,
lissabon	lissabon,lisbon,
australiens	australia's,
nedre	lower,
innanför	inside,within,
minuter	minutes,
vänstra	left,
hästens	horses,horse's,
paraguay	paraguay,
tolkningen	interpretetation,
omloppsbanor	orbits,orbit,
campus	campus,
vinner	gaining,wins,
manlig	male,manly,
identitet	identity,
särskilda	specific,special,
proteinet	protein,the protein,
proteiner	proteins,
illa	bad,
picchu	picchu,
stimulans	stimulating,
betonade	emphasized,
uppfattas	be perceived,are regarded,
försämrades	worsened,worsening,
uppfatta	apprehend,perceive,
sjön	lake,
tämligen	fairly,
astronomi	astronomy,
variation	diversity,
koncentrationsläger	concentration camp,concentration camps; kz-camps,
akademisk	academical,academic,
ärkebiskop	archbishop,
philips	philips,
fakta	facts,fact,
winnerbäck	winnerbäck,winnerback,
baker	baker,
svag	weak,
uppfattningen	comprehension,
framför	above,
förbundet	the union,
okänd	unknown,
nelson	nelson,
mäktiga	powerful,
nederländerna	the netherlands,
båt	boat,
resor	travels,
påsk	easter,
arkitekt	architect,
antisemitiska	antisemetic,anti-semitic,antisemitic,
ozzy	ozzy,
granskning	review,
anfallet	the attack,attack,
huvudstad	capital city,
paris	paris,
tillväxten	growth,
kapacitet	the capacity,capacity,
under	during,under,
läge	location,
svårare	harder,
nordost	north east,the northeast,
pommern	pomerania,
ägande	owning,ownership,
jack	jack,
invånare	resident (-s),inhabitants,
evert	evert,
myntade	coined,
tagit	taken,received,
school	school,
utmärks	are characterized,characterized,
utmärkt	excellent; superb; marked by; characterized by,
öppna	open,
minskar	diminishing,
venus	venus,
matematik	mathematic,
verklig	real,
reklam	advertisement,
parten	party,
markerar	marks,
kropp	body,
bönderna	the farmers,
manus	script,
läget	location,
indierna	the indians,indians,
läger	camps,camp,
stridigheter	oppositions,
aktivt	actively,
drivande	driving,
ebba	die,ebba,
notera	note,
liberty	liberty,
språkliga	linguistic,
aktiva	active,
sund	narrow,sane,
kub	cube,
egyptens	egypts,egypt's,
språken	languages,
zach	zach,
prata	talk,
flera	many,multiple,
medelhavsklimat	mediterranean climate,
utredning	investigation,
beck	beck,
parlamentariska	the parliamentary,
preparat	preparations,compound,
studio	studio,
rysk	russian,
sommartid	summer-time,during summer,
komplex	komplex,
studie	study,
språket	language,
forum	forum,
ty	for,
precis	precisely,exactly; precisely,
svante	svante,
gällande	regarding,
koloniserades	is colonized,colonized,
upptäckter	discoveries,
upptäcktes	discovered,(was) discovered,
julie	julie,
erektion	erection,
övers	translation,
nazistiska	nazi,
misslyckats	failed,
upptäckten	the discovery,
försvarsmakt	armed forces,
eftervärlden	the world,
volym	volume,
klassas	classified,
vinst	profit,win,
miniatyr|px|en	miniature,
konserterna	the concerts,
västtyskland	västttyskland,west germany,
skicka	send,
behandlingar	treatments,
belägg	evidence,
återstående	remaining,
muse	muse,
övertala	convince,persuade,
ludvig	ludvig,
ansökte	applied,
världsarv	world heritage,
fermentering	fermentation,
rörelse	movement,
belgiens	belgium's,
igelkottens	hedgehog,
henri	henri - it's a name,henri,
mm	millimeter,etc.,
arméns	army's,
lukas	luke,
antiken	the ancient world,
ms	motor ship,
mr	herr,mr,
johanssons	johanssons,
avstå	desist,
utgick	started,was deleted,
partiets	the party's,parties,
sträckan	the distance,
utlöste	triggered,
persien	persia,
trädgård	garden,
djur	animals,
genomfördes	was carried out,
fröken	miss,
ena	one,
smält	melted,
iiis	iii's,3's,
väpnade	armed,
ens	even,one's,
gata	street,
elektriskt	electric,
beskrev	depicted,described,
målen	goals,
förståelse	understanding,
mest	mostly,
västvärlden	western world,
målet	the target,
miniatyr|px|ett	miniature,
elektriska	electrical,
frågade	asked,
 cm	centimeters,cm,
nagasaki	nagasaki,
kategorier	categories,
kubanska	cuban,
kontrollen	control,the control,
existera	exist,
arbetat	worked,
arbetar	work,works,
kejsare	emperor,
kampen	the struggle,the fight,fight,
arresterades	was arrested,
vitt	widely,
besittningar	holdings,
synonymt	synonymous,
frivillig	optional,
expansion	expansion,
bibelns	the bibel's,the bible's,
brinner	on fire,burn,
evans	evans,
edith	edith,
nytt	new,
dött	died,
blott	merely,mere,
produktion	production,
upptagen	included,busy,occupied,
livstid	lifetime,
ansvarar	responsible,
alex	alex,
jämförelser	comparison,
detroit	detroit,
bunny	bunny,
ställdes	was positioned,
newport	newport,
storlek	size,
ursprungligen	originally,
erhållit	acquired,received,
önskemål	desire,requests,demands,
gymnasium	high school,
bra	good,
dessförinnan	before (that),before,
träffade	met,
innehållande	containing,including,
platina	platinum,
näst	second,second (to),
nio	nine,
medelålder	middle age,mean age,
behövs	is needed,
kuwait	kuwait,
receptorer	receptors,
användningen	the use,
ammoniak	ammonia,
hemland	homeland,
riktning	direction,
danmarks	denmark's,
paulus	paulus,
behöva	need,
independence	independence,
bröderna	the brothers,
icke	non,none,
fred	peace,
statsöverhuvud	head of state,
samlade	collected,
inom	within,
statsministern	the prime minister,head of state,
studera	study,
tolerans	tolerance,
bredvid	beside,next to,
vetenskapliga	scientific,
samhälle	society,
befolkade	inhabitated,populated,
vetenskapligt	scientifically,
transporterar	carrying,transports,
transporteras	is transported,transported,
nyheter	news,
säsong	season,
museet	the museum,
museer	museums,
föreslagits	was suggested,
nhl	nhl,
institutioner	institutions,
rikaste	the richest,richest,
tillåts	is allowed,allowed,
återvände	returned,
sexuella	sexual,
tillåta	allow,
vikingar	vikings,
tor	thor,
yngste	youngest,
punkten	the point,
à	river,
konventionen	convention,
merkurius	mercury,
å	river,of the,
konventioner	conventions,
ton	tone,
punkter	points,
tom	tom,
uppkommit	arisen,
tog	took,
flertalet	majority; plurality,several,
ifrågasatts	is questioned,
livealbum	live album,
skildes	separated,
meddelande	message,
rädsla	fear,
fördel	advantage,
infaller	falls,
territoriella	territorial,
dramer	plays,
slutsats	conclusion,
mjölk	milk,
uppmuntrade	encouragement,
rad	range,line,
nedgång	decline,fall,
flyttades	moved,
tänka	think,
rak	linear,
somliga	some people,some,
störningar	interruptions,disorder,disorders,
växer	grows,
ras	race,
adhd	adhd,
övervikt	obesity,overweight,
motståndaren	the opponent,adversary,
industriellt	industrial,
hittats	found,
kvällen	the evening,
situationer	situations,
lanseringen	the release,launch,
viktor	viktor,
fartyg	ship; vessel,ship,
industriella	industrial,
planeterna	the planets,the planet's,
mekaniska	mechanical,
grundskolan	elementary school,
tvingas	forced,
skepp	ship,
elektricitet	electricity,
fralagen	fra law,the fra law,
motsatt	opposite,
framgångsrik	successful,
tanzania	tanzania,
sekt	sect,
metan	methane,
sjöar	lakes,
inflytande	influence,
rikskansler	chancellor,
agnes	agnes,
utkanten	the outskirts,outskirts,
dyrare	more expensive,
idrott	sport,sports,
saga	saga,
järnvägarna	the railways,
queen	drottning,
gränserna	borders,the borders,
radio	radio,
höjdpunkt	highlight,climax,high point,
sagt	said,i have said,
radie	radius,
absolut	absolute,
turkar	turks,
claude	claude,
florens	florence,florens,
vinna	win,
ägare	owner,
gods	domain,
holländska	dutch,
abu	abu,
återstår	remains,remain,
andras	others,
länder	countries,
torah	torah,
kommunisterna	communist,the communists,
guatemala	guatemala,
gogh	gogh,
haiti	haiti,
europaparlamentet	european-parliament,the european parliament,
ålder	age,
stadskärnan	town/city,city bear man,
taubes	taubes,
ändras	be changed,
ändrar	changing,changes,
ursäkt	excuse,
ändrat	changed,
lovat	promised,
publicerades	published,
tidningen	the newspaper,paper,
utvisning	penalty,
kroppen	body,the body,
sakta	slowly,
ockuperat	occupied,
fördomar	prejudice,prejudices,
kristendomen	chritianity,christianity,
utformade	designed,
behålla	keep,
mur	wall,
indoeuropeiska	indo-european,european,
brinnande	burning,
antikens	the ancient's,ancient,
populär	popular,
slottet	castle,the castle,
finger	finger,
allra	very,most,-most; most,
mun	mouth,
förhållande	(in) comparison (to),
seder	custom,
betonar	stress,emphasize,
maniska	manic,maniac,
seden	the seed,custom,
dödsorsaken	cause of death,
nummer	number,
kreativitet	creativity,
autonomi	autonomy,
anfall	attack,
verka	seem,operate,appear,
lösningsmedel	solvent,
läggs	put before; submitted; put,lay,
farliga	dangerous,
allierades	allied's,
begränsade	limiting,
förbränning	combustion,
avgöra	determine,decide,
lägga	lay,
grupper	groups,
hitler	hitler,
solljus	sun light,sunlight,
skapades	generated,created,
rumänien	romania,
reglera	expell,controlling,
möjliggjorde	made possible,allowed,
hastighet	speed,
diktatorn	the dictator,
homosexuell	homosexual,
skalan	scale,
öster	east,
modernare	mor modern,
anspråk	claims,claim,
spritt	spread,
drömmar	dreams,
invasionen	the invasion,
älgen	elk; moose,
petrus	petrus,
depp	depp,
förståelsen	the understanding,
nationer	nations,
född	born,
darwins	darwins,
därigenom	by which,thereby,
vojvodskap	voivodeship,
brott	crimes,crime,
maya	maya,
känsliga	1st&2nd: fragile 3rd: sensitive,
nationen	the nation,
kartan	the map,
vanföreställningar	delusions,
varefter	whereafter,
ekonomin	economy,
väljs	elect,
äger	owns,
pekar	points,pointing,
växter	plants,
ökade	increased,
ersatte	replaced,
pekat	pointed,
negativ	negative,
welsh	welsh,
hundra	hundred,one hundred,
formatet	the format,size,
ersatts	replaced,(has been) replaced,
yngsta	youngest,
återvända	return,
uppsving	boost,
gudom	deity,
dylan	dylan,
charlie	charlie,
spelad	played,
svavel	sulphur,
kemikalier	chemicals,
fattigare	poorer,
louisiana	louisiana,
jean	jean,
spelat	played,
spelas	played,
mytologin	mythology,
kraftigt	heavily,
järn	iron,
mängd	volume,
graden	the degree,degree,
sträckor	distances,
grader	degrees,
utföras	performed,
kolväten	hydrocarbons,the hydrocarbon,
kalifornien	california,
använt	used,
värnpliktiga	conscripted,
gavs	gave,
eld	fire,
grundaren	the founder,founder,
aktiv	active,
rätta	correct,come to grips; court; correct,
regionerna	regions,
enlighet	according (to),according,
benämning	term,
donau	the danube,donau,
ämnet	subject,
tillgänglig	available,
kristi	christ,
auktoritet	authority,
ämnen	substances,
gift	married,
såväl	both,as well as,
ladda	load,
modersmål	native language,mother tongue,
bosnienhercegovina	bosnia-hercegovina,
specifik	specific,
tillåtna	allowed,
fotbollen	soccer,
hund	dog,
gifter	marries,toxins,
lagstiftningen	law-making,legislation,
varianterna	the diversities,
hanhon	he/she,
hushåll	household,
besöka	visit,
jennifer	jennifer,
malaysia	malaysia,
besökt	visited,
saturnus	saturnus,
motsatsen	the opposite,
estetik	esthetics,
ultraviolett	ultraviolet,
totalt	complete,wholly,
användare	users,
diktatur	dictator,dictatorship,
utse	appoint,name,
totala	total,
karaktäriseras	characterizes,is characterised,is charactarized,
elitserien	elite series,elitserien,
monoteism	monotheism,
ishockeyspelare	ice hockey player,hockey players,
tillbringar	spends,
män	men,
spelare	player,
hotellet	the hotel,
meyer	meyer,
census	census,
titeln	the title,title,
tvingades	forced,
systrar	sisters,
omgången	round,
plus	plus,
internationell	international,
tydliga	obvious,
genomslag	breakthrough,
primitiva	primitive,
civil	civil,civilian,
menade	meant,
systemet	the system,
tydligt	clear,obvious,
isberg	ice berg,iceberg,
sinne	mind,
anorexia	anorexia,
oförmåga	inability,
omges	surrounded,
omger	surrounds,surrounding,
lagt	laid,added,
kjell	kjell,
sicilien	sicily,
anderson	anderson,
kronprinsessan	crown princess,
metabolism	metabolism,
wittenberg	wittenberg,
föreställa	imagine,pretend; imagine,
fadern	the father,
skulden	the debt,the guilt,
barrett	barett,
fängelsestraff	imprisonment,
italien	italy,
skulder	debts,debt,
finns	is,exist,there is,
fusionen	the fusion,
säkerhet	safety; security,security,
amerikanerna	the americans,
värvade	recruited,
tillika	also,
araber	arabs,
regler	rules,
bildt	bildt,
prov	test,
everest	everest,
bilda	form,
hamn	harbour,
tronen	the throne,
kambodja	cambodians,
förbud	prohibition,
liberalism	liberalism,
tätorten	conurbation,
ni	you,
tillverkade	manufactured,made,
tim	tim,
tio	ten,
lösas	solved,
nr	no.,number,
tätorter	urban,conurbation,cities,
nu	now,
phoenix	phoenix,
sätts	turned (on),is placed,
korrekt	correct,
gäster	guests,
tunna	thin,
massakern	massacre,
cooper	cooper,
kronprins	crown prince,
väckte	awakened,aroused,
beroendeframkallande	addictive,
vietnam	vietnam,
cellens	the cell's,cell's,the cells,
rom	rome,rom,
ron	ron,
rob	rob,
uppskattar	estimates,
rod	rod,
dvärg	dwarf,
knutsson	knutsson,
koreanska	korean,
udda	odd,
minska	reduce,
laura	laura,
mottagarens	the reciever,the receivers,the receiver's,
konstitutionell	constitutional,
bär	berries,here,
tanke	in light of,
federation	federation,
även	even,also,
läns	county's,
varvid	in which,
underhållning	entertainment,
vladimir	vladimir,
krossa	crush,
metod	method,
inlärning	learning,
brother	brother,
olyckor	accidents,
lever	living,live,
der	german word,
försvara	research be,defend,
införandet	the introduction,
trend	trend,
stilar	styles,
kategorirock	category:rock,category rock,
colin	colin,
svartån	svartån (black stream),svartån,
förorter	suburbs,
port	gate,
uppgifterna	the information,data,
ifråga	in question,
poesi	poetry,
agnosticism	agnosticism,
miniatyr	miniature,
ögat	eye,
dem	those,
månaderna	months,
angelina	angelina,
gräs	grass,
kamp	struggle,fight,
vindkraftverk	wind power station,wind turbine,
enkla	simple,single,
utifrån	from the outside,from,
eiffeltornet	the eiffel tower,
jord	soil,
turister	tourists,
dublin	dublin,
införts	introduced,
vägg	wall,
ankomst	arrival,
tilltagande	increasing,
rafael	rafel,
luften	air,
sikt	run,
trummor	drums,
bolaget	the company,
ungerska	hungarian,
russell	russell,
undan	away (from),
utropades	proclaimed,was proclaimed,
samfundet	the communion,
lp	lp,
anda	spirit,
inblandade	involved,
andy	andy,
kurder	kurds,
australian	australian,
turné	tour,
crüe	crüe,
uppskattningar	estimates,
typerna	the types,types,
kär	in love,
övergå	transition,transend,
palestinsk	palestinian,
årets	the year's,
efterhand	hindsight,
piano	piano,
styras	guided,steered,
stater	states,
läkemedel	medicine,
musikaliska	musical,
rådgivare	counsellor,advisor,
valla	valla,herd,
jude	jew,
allvarlig	serious,
domkyrka	cathedral,abbey,
humle	hop,
generell	general,
karibiska	caribbean,
musikaliskt	musically talented,musical,
springsteens	springsteen's,springsteens,
uppväxt	growing up,
bönorna	beans,
dokumenterade	documented,
utdelades	distributed,
hemligt	secret,
annorlunda	different,
hemliga	secret,
ansågs	seemed,
frivilligt	voluntarily,voluntary,
speglar	mirrors,
avrättning	execution,
frivilliga	voluntary,
andlig	spirtual,
stöter	thrust,
simning	swimming,
regeln	the rule,rule,
muslimerna	muslims,the muslims,
inriktad	focused on,intent,
tvserien	tv series,the tv show,television program,
fascism	fascism,
sydliga	southern,
familjens	the familys,family,
flög	flew,
fenomen	phenomenon,phenomenazaqq,
utrikespolitiska	foreign policy,foreign political,
väntan	waiting,
marknad	market,
kroniska	chronic,
stridande	fighting,warring,
japanska	japanese,
väntat	expected,
väntar	waiting,expect,
faser	phases,
kartor	maps,
bushs	bush's,
orten	the suburb,
födelse	birth,
komplicerat	complicated,
iberiska	iberian,
fasen	phase,
rapport	report,
böcker	useful downloads archive,books,
välja	select,
wallace	wallace,
undervisningen	the education,
klasser	classes,
behandlingen	the treatment,the treament,
spelarna	players,
försvaret	the defense,
marleys	marley's,
passar	suits,
hergé	herge,
femte	fifth,
hamilton	hamilton,
karlsson	karlsson,
tredjedel	a third,
hotar	threatens,
opera	opera,
snabb	instant,
namn	name,
futharkens	futhark,the futhark's,
viggo	viggo,
alternativ	alternative,
hotad	threatened,
färger	colors,
bildning	education,learning,
semifinal	semifinals,semi finals,
förhandlingarna	the negotiations,negotiations,
stående	standing,
valuta	currency,
hoppade	jumped,
amerikansk	american,
åsikt	opinion,
tillhörighet	belonging,belonging; affiliation,
behandlas	treated,
upprepade	repeated,
stortorget	stortorget,the main square,
årliga	annual,
profil	profile,
accepterar	accepts,accept,
accepterat	accepted,
kent	kent,
variant	variant,type,variety,
juldagen	christmas day,
zuckerberg	zuckerberg,
etanol	ethanol,
nått	reached,
hjalmar	hjalmar,
gallien	gaul,
soundtrack	soundtrack,
arbetet	work,the work,
traditionen	the tradition,
motion	motion,
traditioner	traditions,the traditions,
place	place,
någonsin	ever,
politiken	the politics,
hemsida	website,homepage,
begår	commits,
såldes	sold,
självbiografi	selfbiografi,
centralamerika	central america,
george	george,
respekt	respect,
given	given,
ian	ian,
vågor	waves,
skjuten	shot,
bahamas	bahamas,
skjuter	shoots,extend,
givet	granted,
folkmängden	population,
personlighetsstörningar	personality disorders,
spelats	played,
webbplatser	webbsites,websites,
gia	gia,
användandet	usage,
grund	in the context: "på grund" = because of,
montenegro	montenergo,
alan	alan,
kallade	called,
nobelkommittén	the nobel commitee,
hur	how,
hus	house,a house,
webbplatsen	webpage,the website,
population	population,
smeknamn	nickname,
modellen	the model,
balans	balance,
marinen	navy,
löfte	promise,
kontroll	control,
framställning	production,
modeller	models,
bildades	founded,was formed,
hjärtat	heart,the heart,
rena	pure,
mottagare	recipient,receiver,
afrikanska	african,
tiotusentals	tens of thousands,
kromosomerna	chromosomes,the chromosomes,
maten	the food,
rent	true,
jordskorpan	earth's crust,earth crust,the earth's crust,
världen	the world,
avstånd	distance,
förste	chief,the first,
första	first,
ideal	ideals,ideal,
förhållandena	conditions,the conditions,
gustavs	gustavs,
konsert	concert,
periodvis	periodically,
stjärnornas	the star's,
knutna	tied,
fci	fci,
falla	fall,
fria	free,
invånarna	inhabitants,inhabitatants; citizens',
staterna	states,
täckt	covered,
täcks	covered,covers,
lisbet	lisbet,
elektromagnetisk	electromagnetic,
betydande	important,
stövare	beagle,hound,
herren	the lord,
tron	faith,
ronaldinho	ronaldinho,
mänskligheten	humanity,
isolering	isolation,
tros	belived,believed,
tror	believe,think,
bandets	the bands,
berättelsen	story,the story,
tvprogram	tv program,tv-show,
guld	gold,
tidningarna	papers,
flydde	fled,
motivet	the motive,
ovanligt	unusual,rare,
iväg	away,
ovanliga	unusual,rare,
analys	analysis,
berättelser	tales,
webbkällor	websources,webbkällor,web sources,
larsson	larsson,
blommor	flowers,
grundandet	founding (of),
tränaren	the coach,
jazz	jazz,
administrativ	administrative,
nedåt	down; downwards,
väder	weather,
anlände	arrived,
forsberg	forsberg,
mörkt	dark,
tränade	trained,
dramat	the drama,
joker	joker,
republika	republic,
osäkert	uncertain,
baltikum	the baltics,
satte	put,put together,
minnen	memories,
underlätta	ease,facilitate,
kraftigare	more powerfully,
inspelningen	recording,
uppdraget	task; assignment,
tekniskt	technical,
stanley	stanley,
minnet	the memory,
älg	moose,
freden	peace,
fredspriset	peace prize,
utbud	availibility,supply,
skett	happened,
önskade	desired,wished,
översättning	translation,
återigen	once again,yet again,
intresserad	interested,
hämtat	collected,downloaded,taken,
konstnären	the artist,artist,
mellan	between,
antagligen	presumably,
konstnärer	artists,
bekämpa	prevent,combat; fight,fight,
ruiner	ruins,
dödade	killed,
myter	myths,
summa	sum,
sydeuropa	south europe,southern europe,
region	region,
ordagrant	literally,literal,
spindlar	spiders,
lenins	lenin's,
introducerades	introduced,
gjorde	did,
gjorda	made,
pakistan	pakistan,
utgåvor	issues,
period	period,
pop	pop,
fransk	french,
werner	werner,
statens	the government's,
utformning	layout,shape,formation,
hävda	claim,
poe	poe,
skånska	scanian dialect,scanian,skånska,
howard	howard,
folken	the peoples,peoples,
strikta	strict,
förekomsten	existence,presence,
dagarna	the days,
musikstil	music style,
folket	the people,
invaderade	invaded,
anderna	andes,the andes,
sändebud	messenger,
andres	andres,other's,
andrew	andrew,
kapitulation	capitulation,
tiger	tiger,silent,
övrig	other,
minister	minister,
kaos	chaos,
hughes	hughes,
användes	was used,used,
riktade	targeted,
mount	mount,
influenser	influences,
cash	cash,
arnold	arnold,
spreds	spread,
fiende	enemy,
grundlagen	constitution,the constitutional law,
synvinkel	perspective,
universums	the universe's,universe's,
pippi	pippi,
nyare	newer,
knyta	tie,
grönland	greenland,
status	status,
producera	produce,
republikens	republic's,
fysiologi	physiology,
protoner	protons,
persons	a person's,persons,person's,
linjerna	routes,the lines,
göring	goring,
producerad	produced,
vatikanstaten	vatican city,the vatican,
relaterade	related,
modet	the fashion,fashion,
medvetna	aware,
kommunistisk	communistic,
pennsylvania	pennsylvania,
breda	wide,
hårdvara	hardwere,
egentliga	real one,
tjänsten	the service,
nordkoreas	north korea's,
medellivslängd	average lifespan,life expectancy,
arkitekten	the architect,
kopplingen	the connection,
lyckan	the happiness,
helsingfors	helsingfors,helsinki,
listorna	the lists of candidates,the lists,
kommentarer	comments,
actress	online,
ekologiska	ecological,
enligt	according (to),according to,
allmän	general,
möte	meeting,
harrison	harrison,
moçambique	mozambique,
leta	search,
utvinns	extracted,
starka	strong,
ny	new,
rose	rose,
regent	ruler,regent,
rosa	pink,rosa,
utbyte	trade,
starkt	strongly,
lett	led (to),
pendeltåg	commuter train,
delstat	state,
feminism	feminism,
riket	kingdom,the land,whole country,
mesta	most,
vampyren	the vampire,
delhi	delhi,
utrikespolitik	foreign affairs,forgein policy,
uppslagsordet	lexical entry; word,entry word,
möts	meet,meets,
majoritet	majority,
vampyrer	vampires,
riken	the kingdoms,kingdoms,
kommentar	comment,
afrikas	africa's,africas,
kennedy	kennedy,
mexikanska	mexican,
tower	tower,
anföll	attacked,
rammstein	rammstein,
verksamheten	the work,
madrid	madrid,
innebära	mean,
gång	time,once,
passera	pass,
latinet	latin,
alkoholer	alcohols,
verksamheter	operations,businesses,activity,
försvarare	defender,
tiders	days',times,time's,
fiktion	fiction,
inspirerades	(was) inspired,
sitta	sit,
stopp	stop,
härledas	derived,
lärda	literate,savants,
buddha	buddha,
legat	layed,
uppbyggnad	construction,structure,
publicerat	published,
willy	willy,
servrar	servers,
geografi	geography,
tyskt	german,
mandelas	mandelas,mandela's,
tyska	german,
tyske	german,
förbindelser	connections,
on	on,
om	for,if,
indianska	red indian,amerindian,native american,
spelet	the game,
of	av,
artiklar	items,
stand	stand,
hindu	hindu,
os	os,
spelen	the games,games,
befäl	command,
koppling	connection,
cambridge	cambridge,
ansträngningar	effort,
tolkning	interpretations,interpretation,
domstol	court,
burton	burton,
befinna	be,
trådlös	wireless,
medlemsstaternas	member state,member states,
valley	valley,
serbien	serbia,
förrän	until,before,
genomfört	carried out,carried through,
jul	christmas,
inriktning	direction,
uppåt	raised,upwards,
ingredienser	the ingredients,ingredients,
koenigsegg	koenigsegg,
manuskript	script,
varning	warning,
ämbetsmän	bailies,
chaplin	chaplin,
kvinnornas	the women's,
taylor	taylor,
felix	felix,
närmast	nearest,closest,
fjorton	fourteen,
liverpool	liverpool,
ökning	increase,
operation	operation,
köpenhamn	copenhagen,
många	many,
mötley	mötley,
utgifter	expenditure,expenses,
babylon	babylonia,babylon,
bredare	wider,
separata	separate,
grupp	group,
ockupation	occupation,
symbol	symbol,
erövring	conquest,
missbruk	addiction,abuse,
vinnaren	winner,the winner,
observatörer	observers,
symtomen	the symptoms,
villkor	condition,
distriktet	district,
barcelona	barcelona,
erfarenhet	experience,
visby	visby,
ali	ali,
alf	alf,
separat	seperate,separate,
ale	ale,
konsekvent	consistent,consistency,
samhällen	communities,societies,
utomliggande	external; ex-territorial,
sakrament	sacrament,
gärning	deed,
uppdrag	job,missions,mission,
persiska	persian,
funktionerna	functions,the functions,
kapitulerade	surrendered,
röstade	voted,
ögonen	eyes,
gary	gary,
påstående	assumption,
cykeln	there are two meanings in the context - cycle and bicycle,
kvar	left,
löper	runs,
färgerna	colors,
liter	liters,
litet	small,
ansluter	connects,connect,
far	father,
fas	phase,
runtom	throughout,
simpsons	simpsons,
fan	devil,
sony	sony,
redaktör	editor,
liten	small,
unionens	the union,european union,the union's,
tjeckiska	czech,
choklad	chocolate,
helvetet	the hell,
list	cunning,
ingående	enter into,in depth,
förtryck	opression,
lisa	lisa,
hitta	make up,come up, find,
grekland	greece,
ted	ted,
istiden	the ice age,
tex	for example,
design	design,
haag	haag,the hague,
what	what,
enklaste	the simplest,
vaginalt	vaginal,
kinesiska	chinese,
version	version,
spelning	gig,
sur	sour,
mördades	murdered,was murdered,
guns	guns,
fäste	attachment,
dottern	the daughter,
upptäcka	detection,discover,
regerade	reigned,
avrättades	was executed,executed,
fjärdedel	fourth,
upptäckt	discovered,
norden	scandinavia; (nordic area; region),the nordic countries,
upptäcks	discoverd,is discovered,
råder	advises,(that) prevails,
soloalbum	solo album,
kärnvapen	nuclear weapons,
tillhörde	was a part of,belonged to,
magnitud	magnitude,
arabemiraten	united arab emirates,uae,the arab emirate,
snus	snuff,
uppkomst	origin,
kategorispelare	category player,
filmerna	the movies,
stöd	support,
dahlén	dahlén,
syfta	aim,refer,
smak	taste,
socialdemokraterna	members of the social democracy,
anarkism	anarchism,anarchy,
succé	success,
kommittén	the committee,committee,
branden	fire,the fire,
förebild	model,role model,
autonom	independent,
gemensamt	in common,
genomsnittliga	average,
israel	israel,
permanenta	permanent,
cellerna	cells,the cells,
akademiens	the academy's,attend,
glas	glass,
hålet	hole; gap,the hole,
floyd	floyd,
glad	happy,
östra	eastern,
naturligt	natural,
investeringar	investments,
godkänt	approved,
decenniet	decade,
decennier	decades,
kryddor	spices,
förhåller	relate,relates,
naturliga	natural,
värt	worth,
division	division,
duett	duet,
bosatt	resident,
huvudort	principal town,
historiskt	historic,historically,historical,
breaking	breaking,
brittisk	british,
satanism	satanism,satanic,
härstamning	origin,descent,
välgörenhet	charity,
indelade	divided into,
rocksångare	rock singer,
skära	carve,
sven	sven,
tagen	taken,
grundämne	element,
fötterna	feet,their feet,the feet,
ångest	anguish,
fötts	born,borned,
atomer	atoms,
regnar	rains,
anarkistiska	anarchistic,anarchist,
praktiska	practical,
bildade	formed,
tsar	tsar,czar,
homosexuella	homosexual,
grande	grand,
greklands	greece's,
människors	people's,
instabil	unstable,
längs	along,
avvisade	rejected,
september	september,
emmanuel	emmanuel,
gudarnas	the gods',god's,
australien	australia,
längd	length,
retoriska	rhetorical,
islam	islam,
lyder	obeys,
rika	rich,
abbey	abbey,
prag	prague,
stephen	stephen,
argentina	argentina,
jämte	next (to),together with,
fenomenet	the phenomenon,
kategorieuropeiska	europe category,
styret	gate,
medborgerliga	civil,
kärna	core,quarks,
postumt	posthumous award,posthumously,
marcus	marcus,
försöken	trials,attempts,the tries,
journalisten	the journalist,
stilen	style,
slidan	the vagina,vagina,
journalister	journalists,
försöker	tries,
principer	principals,
kustlinje	coastline,
ringar	rings,
drycken	beverage,the drink,
betyg	grades,
hawaii	hawaii,
aldrig	never,
mongoliet	mongolia,
ollonet	penis head,the glans,
därvid	thus; thusly; then,therewith,
europas	europe,
väg	way,
kvinna	woman,
vän	friend,
benjamin	benjamin,
poliser	police (-men; -women),police,
ökad	increase,
islamistiska	islamic,
densiteten	density,
beräknades	estimated,
kritiserat	criticized,criticised,
bära	carry,
ökar	increases,
polisen	police,the police,
faller	fall,
fallet	the case,
stavningen	spelling,the spelling,
konsumtionen	the consumtion,consumption,
fallen	cases,
aminosyror	amino acids,
filosofins	the philosophy,
heinz	heinz,
colombia	colombia,
pablo	pablo,
bland	blamd,
story	story,
spred	spread,
lördagen	the saturday,saturday,
misslyckas	fail,fails,
harris	harris,
stort	large,big,
motiveringen	the motivation,
storm	storm,
kristendomens	the christianity's,christianity's,
stora	large,big,
ecuador	ecuador,
sekunder	seconds,second,
mikael	mikael,
gränser	borders,
poster	positions,
serotonin	serotonin,
framtiden	future,the future,
hotet	the threat,the threath,
fattigaste	poorest,
gränsen	the line,border,
besökare	visitors,
siffra	number,
illegala	illegal,
matcherna	the games,games,
direkt	direct,directly,
kina	china,
pjäsen	play,piece,
dans	dance,
guden	the god,
stjärnan	star,the star,
kategorin	category,the category,
klubb	club,
anläggningar	facilities,
kusin	cousin,
tilldelas	assigned,award,
tabell	chart,
omskärelse	circumcision,
slåss	fight,
wilson	wilson,
bedriver	manage,operate,
inriktningar	direction,
dialekt	dialect,brogue,
jämförelsevis	in comparison,comparatively,
judar	jews,
electric	electic,
dagliga	daily,
park	park,
naturvetenskapliga	scientific,
dagligt	daily,
industrialiserade	industrialized,
agnostiker	agnostics,
sånger	songs,
mineral	mineral,
salt	salt,
influensan	the influenza,
sången	the song,
borgmästare	mayor,
statsskick	polity,
kosovo	kosovo,
tjugo	twenty,
ursprungliga	original,
kolonialism	colonialism,
tilly	tilly,
månen	the moon,
tills	until,
beräkningar	calculations,
canaria	canaria,
bidrog	contributed,
moses	moses,
hit	here,
hiv	hiv,
inklusive	including,
vardera	each,
fattiga	poor,
jobbade	worked,
händer	happens,hands,
himmler	himmler,
solsystemet	the solar system,
budapest	budapest,
utvidgade	expanded,
tvkanaler	tv-channels,tv channels,
mediciner	medicines,
avtal	agreement; deal,contract,
tidszon	timezone,time zone,
vincent	vincent,
norrköping	norrköping,
poäng	score,point,
virginia	virginia,
utsatt	exposed,
bars	carried,
etiopien	ethiopia,
art	kind,art,
bart	bart,
arv	heritage,
fiske	fishing,
bara	only,
arg	angry,
stjäla	steal,stealing,
arm	arm,
barn	child,
pär	pär,
bortsett	except,apart,
planeras	is planned,planned,
planerar	is planning,
uppskatta	estimate,appreciate,
inga	no,
planerat	planned,
mördad	murderd,
invaldes	elected,was elected,
planerad	planned,
muslim	muslim,
verksamhet	work,
där	were,
intäkter	incomes,
opposition	opposition,
uppkom	arose,
godkändes	was approved,
tiderna	the times,times, ages,
startades	started,
lyssnar	listen,listens,
roman	novel,
lägret	the camp,camp,
hypotesen	the hypothesis,hypothesis,
lära	get to know,learn,
borta	gone,away,
vidare	moreover,further,
lärt	learned,learnt,
stärktes	was strenghten,
belägna	located,
besegrade	defeated,
östtyskland	east germany,
slott	castle,
hypoteser	hypotheses,hypothesis,
ps	ps,
java	java,
läsa	read,
skrev	said,
personalen	the staff,
kungafamiljen	the royal family,
johannes	johannes,
pc	pc,
byxor	pants,
resultat	result,
ph	ph,
pi	pi,
chandler	chandler,
flight	flight,
togs	taken,were taken,
publiken	the audience,
sydafrikas	of south africa,south africa's,
rättigheterna	the rights,rights,
gården	courtyard; house; farm (-house),
konflikter	conflicts,
konflikten	the conflict,conflict,
deltog	participated,
julius	julius,
sådan	such,kind of,
inspelningar	recordings,
ägs	is owned,(is) owned,
ris	rice,
sjöarna	the lakes,
byggnaderna	buildings,the buildings,
skeppen	the ships,
fysisk	natural,physical,
demografi	demographics,demography,
tidpunkten	the time,the moment,
ideologier	ideologies,
listor	lists,
förföljelse	persecution,
lokal	local,
spears	spears,
låtit	let,ordered,
skeppet	the ship,
byar	villages,
skåne	skåne,scania,
uppbyggd	structered,built-up,
författare	author,
berömt	famous,praised,
kokpunkt	having a boiling point,boiling point,
vinklar	angles,
finansiera	finance,
italiensk	italian,
sjunga	sing,
höjer	rises,raising,
hjärta	heart,
vetenskapen	the science,
kyrkans	the church's,
alfabet	alphabet,
uttalande	statement,
kontinentala	continental,
komplett	complete,
konstitution	constitution,
påverkade	influenced,affected,
remmer	remmer,
dåtidens	past times,that time,
namnet	the name,
folkräkning	head count,
skalv	quake,
minoriteter	minorities,
bostad	lodge,
omedelbar	immediate,
försvunnit	disappeared,
skall	shall,
kongokinshasa	democratic republic of the congo,
minoriteten	minority,
idé	regard,
namnen	the names,names,
skala	scale,scale; size,
färdiga	completed,finished,
synnerhet	specially,particular,
djupare	deeper,
rastafarianerna	the rastafarian,n/a,
begravdes	buried,
användas	used,
stoppade	stopped,
upplevelse	experience,
exakt	precise,
våldsamma	violent,
näringsliv	business,
banbrytande	groundbreaking,
sammansättning	composition,
hittades	was found,
hittas	found,be found,
hittat	found,
minskning	reduction,decrease,
norrut	north,
sjöfart	sea voyage,navigation,
kongo	congo,
lettland	latvia,
trummis	drummer,
global	global,
krigare	warrior,
flottan	the fleet,the navy,
låtarna	the songs,
ungefär	approx.; approximately,approximately,
föräldrar	parents,
grekerna	greek,
statyn	the statue,
frälsning	salvation,
fungera	act,
anne	anne,
trinidad	trinidad,
anna	anna,
höjder	heights,
turism	tourism,
diamant	diamond,
palmes	palme's,plame's,
ställningen	position,
tävlade	competed,
presenteras	was presented,presented,
anklagades	accused,
bayern	bayern,
judendom	judaism,jewism,
kostnaderna	costs,
grundläggande	primary,fundamental,
påtryckningar	pressure,pressures,
tätt	tightly,
vägarna	roads (roadways),
dialog	dialogue,
täta	close,
socialistisk	socialistic,socialist,
oktoberrevolutionen	the october revolution,october revolution,
genomföras	carry out,
medborgarna	the citizens,citizens,
reglerna	rules; regulations,
hållet	way,
abbas	abbas,
km²	square kilometre,
laget	the team,
håller	holds,
dricka	drink,
fast	though; although; fixed; permanent,even though,
jugoslavien	yugoslavia,
bagge	ram,
bruk	use,
ateister	atheists,
delning	division,
rasade	collapsed,
regionen	the region,
längtan	longing,
sköter	handles,
kritikerna	critics,the critics,critiques,
delta	participate,
regioner	regions,
junior	junior,
karolinska	karolinska (institute for medicine),caroline,
anklagelser	accusations,
planeternas	the planets,the planets',
omvärlden	surrounding world,
styrande	rulers,
aktier	stock,
erövrades	conquered,(was) conquered,concoured,
guyana	guyana (name),guyana,
tolka	interpret,
fick	got,was,
z	z,
tidens	time's,that time's,
svenskspråkiga	swedish speaking,swedish-speaking,
ägdes	owned,
singlarna	the singles,
tidpunkt	date,time,
intressanta	interesting,
rainbow	rainbow,
stadion	stadium,the stadium,
liechtenstein	liechtenstein,
psykoterapi	psychotherapy,treatment,
operan	the opera,
mötet	the meeting,
möter	meets,meet,
urval	selection,
skyddas	(is/are) protected,
skyddar	protects,
sutra	sutra,
beräknas	estimated,
beräknar	calculates the,values,
tittarna	the viewers,
stadigt	stable,steadily,
konvertera	convert,
betyder	means,
råkar	happens,happens to,
jugoslaviska	jugoslavian,yugoslavian,
klubbens	club,
oväntat	unexpectedly,unexpected,
underlättar	make it easier,
vice	vice,
europeiska	european,
parallella	parallel,
mesopotamien	mesopotamia,
nasa	nasa,
karma	karma,
lagstiftning	law-making,
nash	' nash,nash,
förhandla	negotiate,
psykologi	psychology,
kanal	channel,
arten	species,
steve	steve,
jimi	jimi,
låter	let,
moseboken	genesis,
norrköpings	norrköpings,
simon	simon,
uppmaning	call; injunction,exhortation,
fortfarande	still,
romerna	the romani,the romani people,
generellt	generally,
generella	overall,general,
hinduism	hinduism,
fotnoter	footnotes,
varierar	varies,vary,
vapen	weapon,
varierat	varied,
sjukdomar	diseases,
medverkade	participated; contributed,participated,
kommitté	committee,
avslutas	close,ends,
avslutat	completed,finished,
tvinga	force,
historikern	historian,the historian,
fiktiva	romantic,
demokratiskt	democratic,
äta	eat,
byggt	built,
noter	notes,
byggs	under construction,
sällsynt	rare,
utanför	outside,
melodier	melodies,
broar	bridges,
demokratiska	democratic,
bygga	build,
indirekt	indirect,
skadad	damaged,
åtminstone	at least,
århundradet	century,
skadan	the hit,the damage,
influerad	influenced,
anderssons	anderssons,andersson's,
skadas	damaged,
västlig	western,
konstant	constant,
folk	people,
influerat	influenced,
hölls	was held,was,
assisterande	assistant,assisted,assisting,
kris	crisis,
skrivna	written,
judy	judy,
krig	war,
dramatiska	dramatic,dramatical,
bröts	was fractured,broke,
koloni	colony,
hdmi	hdmi,
producenten	the producer,
turismen	the tourism,
producenter	producers,
diamanter	diamonds,
filosofi	philosophy,
astrid	astrid,
tvingats	forced,
buddhistiska	buddhistic,
ukraina	ukraine,
metro	metro,
innehar	holds,holding,
innehas	occupied,
innehav	holdings,owning,
anpassat	adapted,
plattan	plate,the plate,
fortsätter	continues,continue,
populärkulturen	popular culture,
egenskaperna	the qualities,
översättningar	translations,
tjänar	serves,
zlatan	zlatan,
reda	find out,find our,
gemenskap	fellowship,
föreställande	depicting,
motor	engine,
redo	ready,
varpå	thereafter,after which,
from	from,
bestämmelser	regulations,
usa	the usa,united states of america,usa,
fel	faults,
fem	five,
sevärdheter	attractions,
upplöstes	dissolved,
källorna	the sources,
inlandet	inland,the inland,
sorg	grief,
andliga	spiritual,
penis	penis,
införande	introduction,
hindrade	preventing,prevented,
vägrade	refused,
fungerar	functions,
reguljära	regular,
beskriva	describe,
automatiskt	automatic,
beskrivs	described,
tar	takes,
tas	is taken,
föreslår	suggest,
ledamöterna	the commissioners,commisioners,the members,
crick	crick,
engels	engels,
tal	speech,
kanadensiska	canadian,
omvänt	reversed,
löften	promises,
beyoncé	beyoncé,beyoncè,
brian	brian,
sig	itself,
sin	its,
väpnad	armed,
kostym	costume,
kontroversiellt	controversial,
roterande	rotating,
oavsett	regardless; whether; irrespective of,regardless,
tack	thanks,
religiös	religious,
bertil	bertil,
lätta	light,lighten,
kontroversiella	controversial,
eritrea	eritrea,
light	light,
centralorter	regional centers,
kommunikationer	communications,
företag	company,companies,
jolie	jolies,
besegrat	defeated,
mekka	mecka,
blandad	mixed,
skapande	creating,creative,
elin	elin,
elit	elite,
blandat	mixed,
karlstad	karlstad,
blandas	mixes,
spotify	spotify,
stiga	rise,
uppmärksammad	noted, come to attention,
förekomst	presence,
befolkning	population,
återvänt	returned,
permanent	permanent,
genomsnittlig	average,
lärjungar	disciple,disciples,
thåström	thastrom,
skede	period,
cypern	cyprus,
betalade	paid,
underjordiska	underground,
fler	more,
östtimor	east timor,
komma	get,
växande	growing,
konungariket	kingdom,
mätt	measured,
studios	the studio's,
boende	resident,housing,
säsonger	seasons,
barnets	the childs,the child's,
byter	changes,exchanges,
kvarteret	quarter,the neighborhood,
säsongen	season,
studion	studio,the studio,
kritik	criticism,critisism,critique; criticism,
alger	algaes,
förbjuda	forbid,ban,
uggla	owl,
minskad	decreased,reduced,
hantverkare	handy worker,craftsman,
från	from,
svar	answer,
bål	torso,
nobelpristagare	nobel laureate (-s); nobel prize winner (-s),
minskat	decreased,
uppnå	achieving,achieve,
plural	plural,
förutsättningar	(pre-)conditions,condition,
hörs	heard,
hört	heard,
hjälpt	helped,
vulkanutbrott	volcanic eruption,
utmärker	characterizes,characterized,
höra	hear,
york	york,
van	van,
philip	philip,
domare	judge,
hörn	corner,
fotbollslandslag	national football team,
gångna	past,past; gone,
tyst	quiet,silent,
waterloo	waterloo,
g	(g),
barns	childrens,children,
via	through,
adrian	adrian,
tvserier	tv-shows,tv shows,tv-series,
tysk	german,
rudolf	rudolf,
ovanpå	on top of,
revolutionens	revolution,the revolutions,
isbn	isbn,
brasilien	brazil,
nietzsches	nietzsche,nietzsche's,
värsta	worst,
regenter	monarchs,
skyddade	protected,
nätverk	network,
enkelt	simple,
åtskilliga	several,
fågelhundar	bird dogs,
meddelanden	messages,
omfattning	extent,
misslyckande	failure,
sankta	sankta,saint,
diskutera	discuss,
rösträtt	right to vote,
valde	crowned,chose,
valda	chosen,
academy	academy,
juli	july,
vind	wind,
dödligheten	mortality,
resterande	remaining,
franska	french,
holland	holland,
franske	the french,french,
birgitta	birgitta,
tommy	tommy,
framgång	success,
algeriet	algeria,
franskt	french,
tomma	empty,
tyskarna	the germans,the german,
heydrich	heydrich,
romarna	the roman,the romans,
cohen	cohen - it's a name,cohen,
benny	benny,
avgörs	determined,is determined,decided,
blir	become,is,
gäng	group,
intervju	interview,
storbritannien	great britain,
byggas	built,build,
uppfann	invented,
lopp	course, passage,races,race,
ansåg	thought,
besittning	dominion,
protesterade	protested,
betydligt	significant,
centra	center,
ström	stream,
centre	center,centre,
who	who,
landslaget	the national team,
intogs	was taken,was captured,
representation	representation,
staternas	states,the state's,
öken	desert,
förbundsrepubliken	the federal republic,federal republic,
undersökte	investigated,examined,
regeringschef	head of government,
miljontals	millions,
enbart	only,
generna	the genes,
moberg	moberg,
uefa	uefa,
blandade	mixed,
funktionella	functional,
debatt	debate,
julafton	chistmas eve,christmas eve,
pastoral	pastoral,
komplicerad	complicated,
dödades	killed,
filmen	the movie,
rösten	voice,the voice,
filmer	movies,
röster	votes,
beroende	dependent,dependent on,depending,
hållning	attitude,
allmänhet	in general,general,
träffa	meet,
gränsar	borders (to),
heta	hot,be named; be called,be called,
överens	in agreement,agree,
gudar	gods,
linje	line,
presley	presley,
hett	hot,
närstående	relative,relatives,kindred,
samtycke	approval,
städer	cities,
mona	mona,
begäran	request,
förbinder	connects,
torka	dry,
mestadels	most of the time,mostly,
kvinnorna	the women,women,
berömd	famous,
nationernas	the nation's,the nations,
rikare	richer,
motståndare	opponents,
theta	theta,
funktion	function,
upplysning	the enlightenment,
praktisk	practical,
sydstaterna	the southern states,southern united states,
vandrar	wanders,migrates,
joe	joe,
swift	swift,
jon	jon,
sångaren	the singer,
allsvenskan	headlines,allsvenskan,
påtagligt	substantially,considerably,
utvecklingen	development,the development,
teoretiker	theorists,
kolhydrater	carbons,carbohydrates,
april	april,
västerländsk	western,
brons	bronze,
vattnets	the water's,the waters,
bronx	bronx,the bronx,
organisation	organization,
betecknar	represent,denotes,
betecknas	designate,labelled,denote,
kategorityska	category: german,
exakta	exact,
korruption	corruption,
vittne	witness,
publicerad	published,
walt	walt,
cirka	approximately,
styrkor	strenghts,forces,
publiceras	publishes,will be published,
framträdanden	appearances,
kuriosa	bric-a-brac,trivia,
utkom	issued,(was) issued,published,
klara	clear,
dödshjälp	euthanasy,euthanasia,
nåddes	reached,
kopplade	connected,
bbc	bbc,
beskrivning	description,
månar	moons,
marilyn	marilyn,
klart	finished,done,
månad	month,
strindbergs	strindberg's,
ständig	constant,
naturtillgångar	natural resources,
mike	micke,
pengar	money,
nickel	nickel,
klassen	the class,
turneringen	the tournament,
dominera	dominate,
lutherska	lutheran,
försvann	disappeared,
fortsättningen	the continuation,
neutrala	neutral,
deklarerade	declared,
plikter	duties,
godkännande	approval,authorization,
bråk	brawl; fight,fights,
problemen	problems,the problems,
officiell	official,
största	biggest,largest,
anpassa	adjust,adapt,
fördelade	divided,distributed,
yngre	younger,
wild	wild,
madeleine	madeleine,
folktro	popular belief,folklore,
explosionen	the explosion,
uppfattning	understanding,
bekräftade	confirmed,
syftar	refers,seek to,refer,
motiv	motif,
jehovas	jehovas,jehova's,
röra	move,
uppstå	develop,arise,
ramels	ramel's,
varar	lasts,
buddhism	buddhism,
pojkar	boys,
samband	connection,
odlade	grew,
skickade	sent,
gett	given,
annekterade	annexed,
tvister	conflicts,disputes,
mottagande	reception,
övervägande	the predominant,predominant,
romeo	romeo,
romer	romani people,roma,
student	student,
raka	straight,
rätt	right,
misstag	mistake,
klubbar	clubs,
vilar	rests,
banden	the bound,
terrorismen	terrorism,the terrorism,
undersökningar	surveys; investigations,studies,
närma	move closer,
ekosystem	ecosystem,eco system,
övertyga	convince,
bandet	band,
organisationens	the organizations,
hårdrocken	hard rock,
lön	salary,wage; salary,
singeln	single,singeln,
uppkommer	arises,arises; generated,
möjligheten	the possibility,
rachels	rachels,rachel's,
erfarenheter	experience,
högskolor	colleges,
patrik	patrik,
miljöer	environment,environments,
antisemitism	antisemitism,
rocken	the rock,rock,
brutit	cut; break,broken,
mytologiska	mytholigical,mythological,
jarl	earl,jarl,
genombrottet	break-through,breakthrough,
alldeles	altogether,
hoppa	skip,
bell	bell,
sky	sky,
rättsliga	justice,legal,
engelsk	english,
ske	happen,
ska	will,shall,
fyller	turns,play,turn; fill,
sanskrit	sanskrit,
serveras	is served,
psykoser	psychoses,
färgen	the color,
olle	olle,
älska	love,
press	press,
psykosen	the psychosis,
säljs	sold,
georges	georges,
budet	the bid,the commandment,
miami	miami,
djupa	deep,
huruvida	whether,
sälja	sell,
gorbatjov	gorbachev,gotbatjov,
immunförsvar	immune defense,
finansieras	financed,finansed,
djupt	deeply,deep,
säkra	safe,secure,
juni	june,
tjeckoslovakien	czechoslovakia,
handeln	trade; commerce,trade,
bibliska	biblican,
efterfrågan	demand,
gäst	guest,
export	export,
försvinna	disappear,
skandinavien	scandinavia,
högst	highest,
planering	planning,
trianglar	with triangles,traingles,
gammalt	old,
risker	risk,
undviker	avoids,
setts	seen,
personligen	personally,
stieg	stieg,
låten	the song,
sjunker	sinks,
markera	mark,
utsöndras	secrete,exudes,
uppvärmning	heating,warming,
mitt	my,
slut	end,
dateras	dated,
sommarspelen	summer games,
ljung	heather,
låna	borrow,
pressfrihetsindex	pressfrihetsindex,
substantiv	noun,
tillräcklig	sufficient,enough,
överlevde	survived,
bestämma	decide,
oberoende	independent,
avsnittet	section,episode,
mellanöstern	the middle east,middle east,
saker	things,
reaktionerna	the reactions,reactions,
mäta	compare,
own	egen,
främre	front,
egna	own,custom,
floder	rivers,
någorlunda	fairly,somewhat,
avrättade	executed,
tillbringade	spent,
mäts	is measured,
floden	river,the river,
vidta	take,
flyger	flying,
folkpartiet	peoples party,
konstruktion	construction,
födelsetal	birthrate,birth rate,
flamländska	flemish,
val	choice,elections,election,
upprättas	established,establish,
vad	what,
smeknamnet	nickname,
mäter	measuring,measure,
regisserad	directed,produced,
nordamerikanska	north american,
lundell	lundell,
identifierade	identified,
granne	neighbour,
hundratal	100,hundred,
ingått	been part of,entered,
krigsslutet	end of war; war's end,
stadens	the town's,the citys,city's,
karta	map,
rybak	rybak,
tema	theme,
missnöjet	grievance,discontent,
jenny	jenny,
reaktorn	the reactor,reactor,
problemet	problem,the problem,
stormakter	great power,superpowers,
eu	eu,
utöva	utÖva,exercise,
runor	runes,
året	the year,
illinois	illinois,
rike	kingdom,
normal	normal,
ursprunget	origin,the origin,
åren	the years,years,
intresse	interest,
serbiska	serbian,
behandlar	treats,treat,
tolkas	interpret,
tolkar	views,
shakespeares	shakespeare's,
tvfilm	tv-movie,
mankell	mankell,
taube	taube,
ställningar	positions,standings,
markant	considerably,marked,
risken	risk,
nödvändigtvis	by necessity,necessarily,
knappast	hardly,
inledning	introduction,the beginning,
bysantinska	byzantine,
tidning	newspaper,
