vanligast	most,most usual,most common,
nordisk	nordic,
uppemot	almost,up,
stammarna	tribes,strains,
arternas	the species,species,
jihad	johad,
elva	eleven,
invandrare	immigrants,immigrant,
hållas	be,be held,
albumet	album,
slå	beat,hit,
albumen	the albums,
hermann	hermann,
lord	lord,
vann	won,
lyckats	succeeded,
dela	divide,dividing,
syrgas	oxygen,
regional	regional,
upptar	occupies,
portugals	portugal,
skicklig	skillful,
statlig	state,government,
medelhavet	mediterranean sea,mediterranean,
andre	other,
helsingborg	helsingborg,
haber	haber,
befogenheter	authorities,powers,
triangelns	triangle,
urskilja	discern,
sture	sture,
sammansatta	composed,
ungerns	hungary,hungrarys,
hanar	males,
upprätthåller	maintains,maintaining,
åsikten	the opinion,view,
åsikter	opinions,
breddgraden	latitude,parallel,
koffein	caffeine,caffein,
filosofer	philosophers,
aten	athens,
hårda	hard,
biografi	biography,
vägrar	refuses,refuse,
filosofen	the philosopher,
motståndsrörelsen	the resistance,resistance,
regnskog	rain forest,rainforest,
baháulláh	bahaullah,bahullah,
föräldrarna	parents,
valrörelsen	election campaign,
bipolär	bipolar,
kids	kids,
demokratier	democracies,
naturen	the nature,
blåser	blowing,
vicepresident	vice president,
robin	robin,
miljarder	billion,billions,
karin	karin,
systematiska	systematical,
unik	unique,
norsk	norwegian,
marino	marino,
hamas	hamas,
systematiskt	systematic,
ansluta	connect,
dna	dna,
sjukdomen	disease,
strikt	strict,
fuktiga	damp,damply,
music	music,
dns	dns,
fuktigt	moist,damp,
pjäs	piece,
musik	music,
befolkningstillväxten	the population growth,the growth of population,
mercurys	mercury's,mercurys,
holm	holm,
politiker	politician,
slutligen	back end,
bulgariska	bulgarian,
temperaturen	temperature,
rasen	the race,
teman	themes,
temperaturer	temperature,
ofta	usually,often,
avancerad	advanced,
vännen	the friend,
köpa	buy,purchasing,
befolkningsutveckling	population development,population growth,
vågen	the wave,scale,
stommen	body,the foundation,
köpt	purchased,
passagerare	passengers,passenger,
kapitalismen	capitalism,
absoluta	absolute,
vänner	friends,
igelkottar	hedgehogs,
hon	she,
kallare	colder,
hov	court,
how	how,
hot	hot,
pågick	lasted,
folkmusik	folk music,
typen	the type,type,
fylla	fill,
inrikes	domestic,
barbro	barbro,
sedd	seen,
objekt	object,
turkiet	turkey,
sankt	st.,sankt,
typer	types,
stormaktstiden	great power period,
grekiska	greek,
arbeten	works,
deutsche	deutsche,
hemlandet	the home country,the homeland,
wind	wind,
vart	each,
varv	revolutions,dockyard,
ormar	snakes,
vars	whose,
dalí	dali,
organismen	the organism,organism,
vare	either,
varg	wolf,
organismer	organism,
vara	be,
barnet	child,
mabel	mabel,
varm	hot,warm,
publicerade	published,
wales	wales,
målade	painted,
assyriska	assyrian,
fil	master of,file,
avgå	resign,
väte	hydrogen,
hemlighet	secretly,
säljande	selling,
hänga	hang,
närliggande	adjacent,nearby,
silver	silver,
utvecklat	developed,evolved,
utlänningar	foreigners,
utvecklar	develops,
utvecklas	development,
terrorister	terrorists,
tingslag	things type,
debut	debut,
utveckling	development,
tillgängligt	available,
utvecklad	developed,
ingrid	ingrid,
tillgängliga	available,
talade	spoke,
angola	angola,
serier	comics,series,
allan	allan,
utvecklandet	development,
serien	the series,
truman	truman,
axelmakterna	axis,
varken	either,
george	george,
slovenien	slovenia,
försökt	tried,
förändringar	changes,
foundation	foundation,
debatter	debates,
ian	ian,
anarkister	anarchists,
metallica	metallica,
ägnade	dedicated,
sannolikt	probably,probable,
att	that,
sysselsätter	employs,
atp	atp,
skjuten	shot,
malmös	malmö's,malmö,
sydost	southeast,
givetvis	course,naturally,
grannlandet	neighboring,the neighbouring country,
östberg	Östberg,ostberg,
tecknade	drew,
övre	top,
djurgården	djurgården,zoo,
förespråkar	advocate,advocates,
xis	the eleventh's,
master	masters,master,
vågade	dared,
ära	honor,glory,
bitter	bitter,
förändringarna	change,
senaten	senate,
bokstäverna	the letters,letters,
förmögenhet	fortune,wealth,
placerade	placed,
nirvana	nirvana,
påverkad	influenced,affected,
ahmed	ahmed,
skatter	taxes,
upphov	origin,source,rise,
tyckte	found,
påverkan	impact,influence,
tree	tree,
gator	streets,
nations	nation,nations,
påverkat	influenced,affected,
varje	each,
utformningen	the layout,
påverkas	affected,
tretton	thirteen,
obligatorisk	obligatory,mandatory,
försörja	support,
densitet	density,
assistent	assistant,
kriterierna	criteria,
boston	boston,
dricker	drinking,drinks,
filosofisk	philosophical,philosophic,
joakim	joakim,
trakten	the region,region,area,
fasta	solid,
normalt	normally,
östeuropa	eastern europe,east europe,
skaffa	obtain,gain,
förhärskande	prevailing,
hjälpmedel	aid,means agent,
bedrivs	conducted,
katalonien	catalonia,
konserthus	concert hall,concert,
victoria	victoria,
gallagher	gallagher,
medlemsstaterna	member states,
anteckningar	notes,
bedriva	carry,prosecute,
eftersom	because,
thriller	thriller,
övertog	took over,overtook,
annars	else,
singer	singer,
morgon	tomorrow,
arkitektur	architecture,
öland	oland,öland,
camp	camp,
utmärkande	characteristic,distinguishing,
förlorar	loses,
översatt	translated,
förlorat	lost,
grovt	heavy,rough,
passerade	passed,
singel	single,
tänkte	thought,was going to,
inspelning	recording,
ungar	kids,
verkställande	executive,
anorektiker	anorexic,anorectic,
bandmedlemmar	band members,
konkret	specific,concrete,
pris	price,
teater	theater,
louise	louis,
populärkultur	popular culture,
buss	bus,
than	than,
övergår	surpasses,
sekulär	secular,
bush	bush,
omvända	reverse,
rice	rice,
mottog	received,
lastbilar	truck,
storbritanniens	united kingdom,
tillståndet	state,the state,
rättegången	trial,the trial,
årsdag	anniversary,
upprätta	establish,up,
metoden	the method,
dansk	danish,
plats	place,
bensin	gasoline,
lyssna	listening,listen,
balans	balance,
innebörd	meaning,
spänning	voltage,
hantverk	crafts,
×	x,
kallt	cold,
sköta	operate,
utgåvan	the edition,
uppgift	task,data,
framfördes	were,
genomsnittet	average,the average,
release	release,
kalla	cold,
ovtjarka	caucasian shepherd dog,
blev	became,was,
etik	ethics,
flagga	flag,
skulle	could,would,
skriva	write,
bygger	based,
arlanda	arlanda,
skrivs	written,
hedersdoktor	honorary degree,honorary doctorate,
manson	manson,
förhindra	prevent,
wikipedia	wikipedia,
upphovsrätt	copyright,
sundsvalls	sundsvall,
figur	figure,
sista	last,
siste	last,
österrike	austria,
ringa	call,
rollen	role,the role,
henrik	henrik,
ställning	position,
lanserades	was launched,
tilldelades	awarded,
kommunikation	communication,communications,
världsturné	world tour,
roller	roles,
yttre	outer,
tillämpar	practice,administers,
tillämpas	applied,
huvudet	head,
country	country,
sparta	spartans,sparta,
följas	followed,
pitt	pitt,
edgar	edgar,
nordiska	nordic,
nederlag	defeat,
nordiskt	nordic,
genus	gender,genus,
logik	logic,
summan	sum,the sum,
igelkotten	the hedgehog,
folkmordet	genocide,
armén	the army,
herr	mister,
afrikanska	african,
fra	fra,
union	union,
avgörande	settling,essential,
fri	free,
tiotusentals	tens of thousands,
operationer	operations,
socialistiskt	socialistic,socialist,
årtionde	decade,
fru	mrs.,wife,
arbetslösheten	unemployment,
verktyg	tools,
barndom	childhood,
life	life,
café	cafe,café,
ifrån	off,
ändrade	changed,modified,
arkiv	archives,archive,
närvarande	present,
dave	dave,
kometer	comets,
chile	chile,
övergripande	overall,general,
chili	chili,
parterna	parties,
intag	intake,
slutliga	evenutal,
frankrikes	frances,
castro	castro,
klarade	passed,
organisera	organize,organizing,
kontraktet	the contract,contract,
tintin	tintin,
brister	failures,inabilities,
gärna	readily,
desto	the,ever,
stämma	meeting,
player	player,
tänkare	thinker,
australia	australia,
bristen	lack of,lack,
slag	kinds,type,
madonna	madonna,
tät	compact,sealed,
serbisk	serbian,
tillhandahåller	provides,
vrida	twist,turning,
foton	images,photos,
agnetha	agnetha,
european	european,
materiell	material,
funktionen	the function,
josef	joseph,josef,
topp	top,
värde	value,
emi	emi,
föras	be,be brought,taken to,
synder	sins,
tung	heavy,
zeeland	zealand,zeeland,
kampanj	campaign,
gudinnan	the godess,
grundlag	constitution,
försvarade	defended,
manteln	mantle,
snö	snow,
köra	run,drive,
koloniseringen	colonization,
capitol	capitol,
dödsoffer	casualty,death victim,
biskop	bishop,
krigsmakten	armed forces,
körs	driven,being driven,
birmingham	birmingham,
utrotning	extinction,
valutan	currency,
kommunal	communal,municipal,
döda	dead,
givit	gave,
matteus	matteus,
han	he,
grafit	graphite,
vetenskapsmän	scientist,scientists,
bnp	gdp,
ideal	ideals,
muhammeds	muhammad,
huvud	head,
hette	name was,named,
lunginflammation	pneumonia,
har	is,has,
hat	hatred,
hav	seas,ocean,
präst	priest,
underliggande	underlying,
svensson	svensson,smith,
narkotika	drug,narcotics,
livsstil	lifestyle,
bushs	bush,
melodifestivalen	eurovision song contest,
uppmärksammade	observed,
county	county,
bobby	bobby,
sedlar	bills,
alice	alice,
konsert	concert,
residensstad	city of residence,county seat,
sebastian	sebastian,
ola	ola,
old	old,
företräder	representing,
people	people,
billboard	billboard,
parlamentarisk	parliamentary,
delade	split,
kulmen	culmination,the acme,peak,
fot	foot,
for	for,
varierande	varied,varying,
fox	fox,
angränsande	adjacent,
utser	appoints,
utses	is appointed,
akademi	academy,
idéer	ideas,
myndigheter	authorities,agencies,
annan	another,
neptunus	neptune,
stefan	stefan,
påminner	reminds,out,
hörde	heard,
binder	bind,
olympiska	olympic,
möjligheterna	possibilities,the possibilities,
myndigheten	the authority,authority,
annat	alia,other,
evangelierna	gospels,
army	army,
mynnar	opening,
stjärna	star,
misstänkt	suspect,suspected of,
nixon	nixon,
hänt	suspension,happened,
delvis	partial,partly,partially,
döpte	renamed,
psykiska	mental,
marshall	marshall,
som	as,which,
sol	sun,
lagliga	legal,lawful,
son	son,
psykiskt	psychic,mentally,
fci	fci,
delarna	parts,
artikeln	the article,
hantera	handle,
nova	nova,
säkerhetspolitik	safety policy,security,
joseph	joseph,
 miljoner	millions,millon,
jane	jane,
 mm	millimeter,
happy	happy,
saltkråkan	salt crow,
offer	victims,victim,
öppen	open,
förhållanden	relationships,conditions,
öppet	open,
verde	verde,
tigern	the tiger,
avsevärt	substantially,considerably,
drabbat	affected,
gymnasiet	high school,
drabbar	affect,troubles,
polska	polish,
syften	purpose,
pest	plague,
syftet	purpose,
fansen	fans,
moderna	modern,
föregångare	predecessor,precursor,
konung	king,
lunds	lund,lund's,
låtar	songs,
modernt	modern,
krävde	demanded,
ericsson	ericsson,
elektromagnetisk	electromagnetic,
huvudperson	protagonist,
dotter	daughter,
aristokratin	aristocracy,
protester	protests,
läste	read,
republik	republic,
roll	role,
olja	oil,
reggae	reggae,
avskaffades	was abolished,
bostadsområden	residential,housing,residential areas,
palme	palme,
blått	blue,
vintrarna	the winters,
modell	model,
rolling	rolling,
utbildade	formed,
aragorn	aragorn,
tävling	competition,
sällan	rare,
povel	povel,
laddade	charged,
perioden	period,
kategorifödda	category born,
förtjust	fond,delighted,
trettio	thirty,
time	time,
skatt	tax,
erkände	acknowledged,
oss	us,
ost	cheese,
uppgifter	tasks,data,
stödjer	support,supports,
uppgiften	the task,task,
atombomben	atomic bomb,the nuclear bomb,
stålgemenskapen	steel community,
inkomst	income,
machu	machu,
vet	know,
fängelset	prison,
intresserade	interested,
grön	green,
vem	who,
bosnien	bosnian,bosnia,
musikstilar	music genres,music,
individer	subjects,
choice	choice,
individen	the individual,individual,
framställs	is depicted,prepared,
skillnaderna	the differences,differences,
kompositörer	compositors,
initiativ	initiative,
lägre	lower,
inhemska	native,
myntade	coined,
energin	the energy,
oppositionen	opposition,
årig	year old,minor,
jämnt	even,evenly,
nybildade	newly formed,
scen	stage,
jämna	even,
firandet	the celebration,
måne	moon,
greve	count,earl,
elton	elton,
köp	purchase,
kör	run,
kunskapen	the knowledge,
beskydd	conservation,
axel	axel,
bosatte	settled,
kön	gender,sex,
kunskaper	knowledge,
kusten	the coast,coast,
katter	cat,
berättelsen	the story,
provinserna	provinces,the provinces,
galileo	galileo,
vintertid	winter-time,winter,
budskapet	message,
katten	the cat,
huvudsakliga	main,
studien	study,the study,
genomgående	consistently,through,
hälft	half,
studiet	study,the study,
studier	studies,
love	love,
santa	santa,
publicera	publish,
kommit	come,
presenterade	presented,
canis	canis,
sprids	spreads,
samlat	collected,gathered,
samlar	collect,
positiva	positive,
änglar	angels,
vuxna	adult,
sprida	spread,
judarna	jews,
positivt	positive,
samlag	intercourse,
effektiv	effective,
ställt	taken,put,set,
ställs	is,
dagars	day,days,
hår	hair,
tillträdde	took,
ställe	place,
ställa	make,set,
tabellen	table,
dålig	poor,
grönt	green,
straffet	penalty,
mörker	dark,
kunskap	knowledge,
gröna	green,
phoebe	phoebe,
påvisa	detection,show,
stigande	rising,up,
locka	attract,
missförstånd	misunderstanding,misunderstandings,
locke	locke,
släktskap	kinship,
inkluderade	included,
porträtt	portraits,portrait,
utnyttjade	utilized,
svenskar	swedish,swedes,
milda	mild,
årligen	annually,annual,
skikt	layers,layer,
svenskan	swedish,
storleken	size,
trigonometriska	trigonometric,
européer	europeans,
levande	live,
riksdagen	parliament,the parliament,
gigantiska	gigantic,giant,
kungens	king,the king's,
löpande	running,assembly,
svart	black,
nyligen	recently,
data	data,
epost	e-mail,email,
portugisiska	portuguese,
stress	stress,
natural	natural,
bergarter	rock types,rocks,
undervisning	teaching,education,
påstod	claimed,
ss	ss,
sr	sr,
sv	south west,
vikt	weight,
st	saint,
sk	so called,known,
so	so,
sm	swedish championship,
sa	said,
vika	fold,
se	see,
resulterar	resulting,result,
vintrar	winters,
resulterat	resulted,resulted in,
professorn	professor,
kong	kong,
antingen	either,
allvarligt	serious,severe,
clinton	clinton,
irländsk	ireland,
torg	square,
ingvar	ingvar,
dialekter	dialects,
utsätts	exposed,
jim	jim,
tilldelats	assigned,awarded,
begrepp	term,concept,
ersätts	replaced,
faderns	his father,the father's,
monopol	monopoly,
personlig	personal,
britter	britons,
hos	of,with,
änden	end,
öppnades	were opened,was opened,opened,
musiken	the music,music,
matcher	matches,games,
datorspel	video game,computer game,
nation	nation,
records	records,
matchen	the game,
kategoripersoner	category of persons,
kantoner	cantons,
kravet	requirement,the demand,
musiker	musicians,
atmosfär	atmospheric,
lockar	curls,
förväxlas	confused,mistaken,
sidor	sides,
skivkontrakt	record contract,
dominerar	dominate,dominates,
domineras	dominated,
runstenar	runestones,
dominerat	dominated,
födelsedag	birthday,
prisma	prism,
dynamiska	dynamic,
står	standing,star,
stål	steel,
hinduer	hindu,hindus,
krav	requirement,
kött	meat,
riktigt	real,
ockupationen	occupation,
specifikt	specifically,
sjuka	disease,sick,
avgör	decides,determines,
riktiga	real,
bränder	fires,
internet	internet,
roterar	rotates,
bla	blah,among others,
sfären	spheres,sphere,
garantera	ensure,guarantee,
vård	healthcare,
våra	our,
sålde	sold,
bytt	changed,traded,
byts	changed,replaced,
sålda	sold,
väster	west,
pilatus	pilatus,pilate,
dramaten	dramaten,
byta	change,trade,
föreställning	performance,
fyllt	filled,
pund	pound,
artister	performers,
punk	punk rock,para,
flandern	flanders,
solna	solna,
artisten	the artist,artist,
gordon	gordon,
främst	all,primarily,
huvudstäder	capitals,
givits	given,
jakob	jakob,
hård	hard,
one	one,
slutet	end,
tsunamier	tsunamis,
hårt	hard,
open	open,
ont	bad,
urin	urine,
city	city,
teologi	teology,theology,
skådespelarna	actors,
råolja	crude oil,
intill	beside,adjacent to,adjacent,
sjö	naval,lake,
nästa	next,
williams	williams,
animerade	animated,
vilka	who,which,
tillräckligt	sufficient,
irakiska	iraqi,
tillräckliga	insufficient,sufficient,
svenskarna	the swedes,
provins	province,
dygn	day,
fiskar	fishes,fish,
uppenbarelser	revelations,
berlinmuren	berlin wall,
kamprad	kamprad,
motståndarna	the opponents,opponents,
tankar	tank,thoughts,
sak	thing,substance,
san	san,
sam	co,
generation	generation,
konsekvenser	consequences,
argument	arguments,
församlingar	parishs,assemblies,
say	say,
känslan	feeling,the feeling,sense,
allen	allen,
turner	tournament,
staden	city,the city,
priserna	the prices,
övriga	others,
takt	rate,
styrelsen	the board,board,
zoo	zoo,
jefferson	jefferson,
harald	harald,
övrigt	other,
förändringen	the change,change,
föder	gives birth,
muslimer	muslims,
finlands	finlands,
sekreterare	secretary,
tränare	coach,
mynt	coins,coin,
religionen	the religion,
betyda	mean,
religioner	religions,
forskningen	the science,research,
rådets	council,
kontroversiell	controversial,
driva	operate,run,
förändras	changes,
inledningen	the introduction,
ursprung	root,
fredspriset	peace prize,peace price,
rykte	reputation,
färdig	pre,done,
drivs	driven,run,
salt	salt,
olagligt	illegal,
axl	axl,
beckham	beckham,
ledd	led,
dimensioner	dimensions,
dahléns	dahlen,
sjöss	sea,
antalet	number,the number,
stärkte	strengthened,
slog	hit,
hockey	ice hockey,
caroline	caroline,
carolina	carolina,
beatles	beatles,
kategorimusik	category music,
katoliker	catholics,
inlägg	post,
beatrice	beatrice,
egentliga	actual,
platta	flat,
undersöka	study,research,
rörande	concerning,
spetshundar	tip of dogs,
ländernas	the countries,countries,
artist	artist,
råd	council,
enighet	unity,
översättningen	translation,
roger	roger,
varna	alerting,
sträcka	distance,
monark	monarch,
erbjöds	offered,
dagsläget	present situation,current situation,
översättning	translation,
brännvin	schnaps,aquavit,
snabbare	rapid,faster,
behovet	the need,
up	i[,up,
nederbörden	precipitation,the precipitation,
skärgård	archipelago,
talman	spokesperson,
ordspråk	proverbs,proverb,
enhetlig	uniform,
utgörs	consists of,is,
förvaltning	management,
källa	source,
kritiserade	critisized,criticized,
begränsningar	limitations,
upplever	experiencing,experience,
utgöra	compose,make up,
kilometer	kilometer,kilometers,
revolutionär	revolutionary,
små	small,
amerikanskt	american,
anledningarna	the reasons,
screen	screen,
fynd	findings,
antika	ancient,
amerikanske	american,
awards	awards,
amerikanska	american,
mariette	mariette,
basisten	bassist,basist,the basist,
skönlitteratur	nonfiction,
mans	man's,
nationell	national,
rekord	record,
mani	mania,
tillsätts	added,appoints,
långsammare	slower,
upproret	the upprising,rebellion,
klimat	climate,
hamnade	landed,ended up,
drogs	was pulled,was,
därtill	thereto,
teddy	teddy,
farfar	paternal grandfather,
west	west,
bolag	company,
luft	air,
cupen	the cup,cup,
lidit	sustained,suffered,
lånat	borrowed,
förr	sooner,before,
formen	the form,form,
formel	formula,
sångerska	songstress,singer,
diktaturen	dictatorship,
tillåter	allow,
tillåtet	allowed,
former	forms,
landskapen	landscapes,
samling	concentration,collection,
vojvodina	vojvodina,
starkt	strong,
landskapet	landscape,
värderingar	evaluations,values,
situation	situation,
ive	i've,
aston	aston,
bror	brother,
bron	bridge,the bridge,
tillåtelse	allowed,permission,
sammanfaller	coinciding,coincides,
beteckna	denote,
ohälsa	disorders,
världsbanken	world bank,
ståndpunkt	standpoint,position,
träffat	met,
wilhelm	wilhelm,
otto	otto,
träffas	reached,
oceanen	the ocean,ocean,
ekologi	ecology,
ludwig	lugwig,
nationalparker	national parks,
brändes	burned,burnt,
singapore	singapore,
sägas	is said,said,
lindgrens	lindgren's,lindgrens,
följer	resulting,
förkortning	abbreviation,
senator	senator,
dsmiv	dsm-iv,
personlighetsstörning	personality disorder,
måla	target,
tillfälle	occasion,time,
gestalter	figures,
avser	regard,refers to,
avses	regard,
ifrågasatt	questioned,
iraks	iraq,
gudomliga	divine,
summer	sommar,
förluster	loss,losses,
bokförlaget	bokförlaget,
berättelse	tale,story,
rest	residual,
koncentration	concentration,
spårvagnar	trams,
psykologisk	psychological,
resa	travel,
libyen	libya,
förlusten	loss,
heliga	saints,
sprider	spreads out,spreads,
helige	holy,
isen	the ice,
instrument	intrument,
körberg	körberg,
sänka	lower,
infördes	introduced,
unikt	unique,
heligt	holy,
störst	most,
snart	soon,once,
vinkel	angle,
regim	regimen,regime,
unesco	unesco,
litteraturen	literature,
skadade	wounded,damaged,
stammar	strains,stutters,tribes,
statsreligion	state religion,
framsteg	progress,
tvserie	tv serial,
carl	carl,
tsunami	tsunami,
ekonomier	economies,
stupade	fallen,killed,
intet	nothing,no,
jobbar	work,
nämnas	mentioned,include,
domkyrkan	cathedral,
ursprungsbefolkning	native population,indigenous,
ekman	ekman,
kännedom	known,knowledge,
närheten	near,
björn	bear,
västerås	vasteras,västerås,
institutionerna	institutions,
än	yet,than,
exil	exile,
inkluderar	include,includes,
cannabis	cannabis,
varsin	opposite,
är	is,
katolsk	catholic,
långstrump	longstocking,
jacksons	jackson's,jacksons,jackson,
nivån	level,
medlemsstater	member,member-state,
stone	least,
organisationen	the organization,
ace	ace,
herrlandslag	men's national team,women's national teams,
vissa	some,
populationen	the population,population,
befinner	is,
digerdöden	black death,the black death,
populationer	populations,
lyssnade	listened,
organisationer	organizations,
visst	specific,certain,
billboardlistan	billboard list,bilboardlist,
berger	berger,
upplevelser	experiences,
ronden	round,
berget	mount,the mountain,
nationalencyklopedin	national encyclopedia,the national encyclopedia,
tillägg	addition,appendix,
säkerhetsrådet	security,
partiet	the party,portion,
bryta	break,
partier	portions,parties,
lätt	easy,
het	hot,up to date,
företag	company,companies,business,
striderna	fighting,
förintelsen	holocaust,the genocide,
philadelphia	philadelphia,
evangeliska	evangelical,
söker	seeks out,
hel	full,
hem	back,
hamnen	the harbour,
sover	sleep,
enorm	huge,enormous,
hänvisning	reference,
project	project,
dagen	day,
hells	hells,
bevarat	preserve,preserved,
bevaras	are protected,preserved,
kontroverser	controversies,
språkliga	linguistic,
bevarad	kept,preserved,
åttonde	eighth,
rush	rush,
sällskap	groups,
jamaicas	jamaicas,jamaica's,
kvartsfinalen	quarter finals,quarterfinals,
utmed	along,
vinkeln	the angle,
afrodite	aphrodite,afrodite,
förbundsstat	federal,federal state,
produkt	product,
regimer	regimens,regimes,
krona	crown,
ac	ac,
ab	ab,
brodern	brother,
redovisas	reported,accounted for,
gustafs	gustafs,gustaf's,
am	am,
al	alder,
bronsåldern	bronze age,the bronze age,
as	as,
beordrade	commanded,ordered,
at	at,
av	of,
håll	ways,hold,
väsentligt	substantially,relevant,
testamentet	testament,
vore	were,
federala	federal,
rökning	smoking,
innehåll	content,contents,
svårt	hard,difficult,
belönades	awarded,
isolerad	isolation,
avslöjade	revealed,
såsom	such as,
gifta	marry,married,
värmlands	värmlands,
koppar	copper,
gifte	married,
medverkan	participation,
kvarstod	remained,
kategorisvenskspråkiga	category swedish-speaking,
terra	terra,
medverkat	participated,
värd	host,worth,
terry	terry,
ekonomi	economy,
forntida	ancient,prehistoric,
kommunen	municipality,
skador	damage,
århundradena	centuries,
beteckning	label,
nelson	nelson,
decennierna	decades,
original	original,orignal,
renässans	renaissance,
släppt	released,
släpps	released,
elektron	electron,
halsen	throat,the throat,
anpassning	adjustment,
kammare	chamber,
års	years,
släppa	release,
likartade	similiar,similar,
norr	north,
skogarna	the forests,
number	number,
pojkvän	boyfriend,
ullevi	ullevi,
tv	tv,
romanen	novel,
nederbörd	rainfall,precipitation,
to	to,
mildare	milder,mild,
belägg	evidence,
th	th,
nord	north,
te	tea,
sättas	turn,added,
ta	to,take,
avlägsna	remove,
användes	was used,
arvet	the inheritance,heritage,
telefonen	the telephone,
strand	beach,
utländsk	foregin,foreign,
sant	true,
ensamma	alone,
djurarter	species of animals,animal species,species,
borrelia	borreliosis,
muslimska	muslim,
utsåg	declared,appointed,
sand	sandy,
siffrorna	figures,numbers,
områdets	the area's,area,
harry	harry,
sann	true,
språkbruk	parlance,language,
förmedla	pass,
döttrar	daughters,
påståenden	claims,assertions,
synd	sin,
dödsstraff	death penalty,
utökade	expanded,
vägnät	network,
stöder	supporting,
pass	an,
givaren	the giver,
syns	visible,
stängt	closed,
delen	part,
soldater	soldiers,
islams	islams,islam's,
gjorts	made,done,
hänsyn	light,consideration,
full	full,
gruppen	the group,
själen	the soul,
arkeologiska	archaeological,
grupper	groups,
legend	legend,
motstånd	resistance,opposition,
äventyr	adventures,
traditionella	traditional,conventional,
exklusiv	exclusive,
traditionellt	traditional,
social	social,
action	action,
oftare	more often,more,
varelser	creatures,
medlemskap	membership,
kommunistpartiet	communist party,the communist party,
vid	by,in,
ordinarie	permanent,regular,
vin	wine,
hamnat	ended up,got in to,
juridiskt	judicial,
vis	vis,
kuiperbältet	the kuiper belt,
vit	white,
spelaren	the player,
motsatsen	the opposite,opposite,
biskopen	the bishop,
mors	mother,
petroleum	oil,petroleum,
underordnade	subordinates,
pearl	pearl,
sitter	is,serve,sit,
presenterades	presented,
rhen	rhine,
dödligt	lethal,deadly,
mora	mora,
inslag	impact,elements,
mord	murder,
uppskattad	estimated,
berättade	told,
angående	concerning,reference,
uppskattas	is appreciated,estimated,
uppskattar	estimated,estimates,
schweiz	switzerland,
undergång	doom,destruction,
socialt	socially,social,
inträffade	occurred,happened,
medelklassen	middle class,
science	science,
sociala	social,
morgan	morgan,
kapitalism	capitalism,
studenter	students,
läkaren	the doctor,physician,
samväldet	commonwealth,the commonwealth,
nobelpriset	the nobel prize,
säljas	is sold,sold,
nordvästra	northwest,north western,
skadliga	harmful,deleterious,
huvudstaden	capital,
mellersta	middle,the middle,
states	states,
stater	states,
spansk	spanish,
järnvägsnätet	railroad network,rail,
information	information,
vägnätet	road network,
hugo	hugo,
uppfattade	perceived,
ansetts	considered,regarded,
lejon	lion,
riksdagens	the parliament's,the parliaments,
retorik	rhetoric,
fortsättning	continuation,continued,
hustru	wife,
produktionen	production,the production,
lanka	lanka,
komplext	complex,
anklagade	accused,
pucken	the puck,
komplexa	complex,
utvidgning	enlargement,
hållit	held,maintained,
nationerna	the nations,nations,
blommor	flowers,
trade	esterified,
utgjordes	was,
scott	scott,
kvinnors	women,women's,
aktiviteter	activities,activity,
anställda	employed,
radion	radio,
vietnamkriget	the vietnam war,vietnam war,
känsla	feeling,sense,
alla	all,
högskola	college,
protestanter	protestants,
caesars	caesars,
miljön	environment,the environment,
termen	the term,term,
hounds	hounds,
termer	terms,
allt	all,
alls	all,
få	gain,
van	van,
isaac	isaac,
konstruerade	constructed,
samhällets	society,of society,
berömda	famous,
inleda	initiate,
beräkna	calculate,
producerad	produced,
inledande	initial,
produceras	produced,
producerar	producing,
grekisk	greek,
producerat	produced,
introducerade	introduced,
producerade	produced,
olycka	accident,disaster,
intåg	advent,
budskap	message,
målning	painting,
graviditet	pregnancy,
blodet	the blood,
denne	his,
denna	that,
härrör	derived,
enstaka	occasional,single,
england	england,
populärt	popular,popularly,
sydöst	southeast,
doser	dose,
populära	popular,
blues	blues,
förespråkade	advocated,
kretsen	the order,circuit,
finner	found,finds,
uppfördes	was constructed,built,
återkomst	return,
omröstningen	vote,
kopplad	connected to,connected,
garvey	garvey,
avgick	retired,
norska	norwegian,
uppstått	resulting,arisen,
sammanfattning	summary,
besökte	visited,
kopplat	connected,coupled,
kopplas	connected,coupled,
highway	highway,
medel	middle,medium,
sparken	gets fired,fired,
alltmer	increasingly,more and more,
beethoven	beethoven,
stjärnor	stars,
poeter	poets,
driver	run,drive,
båda	both,
både	both,
kostade	cost,
ålands	Åland island's,aland,
kärnkraft	nuclear power,nuclear,
poeten	the poet,
teknologi	technology,
service	service,
turistmål	tourist attraction,
hjärta	heart,
samlas	together,
målningar	paintings,
skolan	school,
nivåer	levels,
besök	visit,
uppenbarelse	apparition,
principen	the principal,principle,
bidragit	contributed,
relationer	relations,
foten	foot,
skiftande	shifting,
spekulationer	speculations,
såg	see,saw,
gemensamma	common,
avel	breeding,
liknas	compared to,likened,
liknar	similar,
tove	tove,
saint	saint,
sår	wound,
missade	failed,
besläktat	related,
läggas	laid,added,
chefen	head,
tappade	lost,
zeus	zeus,
zeppelin	zeppelin,
moder	mother,
svår	severe,
grace	grace,
obama	obama,
organiseras	organized,
återkom	return,returned,
organiserat	structured,
niklas	niklas,
koncentrerade	concentrated,
marknadsekonomi	market,market economy,
freud	freud,
organiserad	organized,
nikolaj	nikolaj,nicholas,
ägg	eggs,
äga	be,
väljer	select,
inkluderas	include,is included,
statyn	the statue,statue,
generationen	the generation,
inkluderat	including,
ägt	taken,
generationer	generation,generations,
astronomin	astronomy,
visats	shown,demonstrated,
framåt	forward,forth,
varianten	version,variant,
norstedts	norstedt's,collins,
kongokinshasa	democratic republic of the congo,congo kinshasa,
varianter	varieties,diversities,
vinterspelen	winter games,
arabisk	arabic,
edison	edison,
sydostasien	south east asia,southeast asia,
brooklyn	brooklyn,
plan	flat,level,
kombinationer	combinations,
arter	species,
utsattes	subjected,exposed,
cover	cover,
kanalen	the channel,channel,
kanaler	channels,
monarki	monarchy,
arten	species,
kombinationen	the combination,
golf	golf,
gold	gold,
omfattade	included,
falska	false,
presidentens	president,the presidents,
detalj	detail,
karaktär	character,
falskt	false,
framgångar	successes,success,
existensen	existence,
betydelser	values,meanings,
jämföra	compare,
wayne	wayne,
betydelsen	the meaning,significance,
jämfört	compared,
kontor	office,
karakteristiska	characteristic,
genomgick	underwent,
gratis	free,
evolutionen	evolution,the evolution,
tekniken	techinque,art,the technology,
tekniker	technician,
actress	actress,
utbildningen	education,
föll	fell,
erkännande	recognition,
victoriasjön	victoria lake,lake victoria,
tanken	the thought,idea,
ledare	conductors,leader,
cry	cry,
populärmusik	popular music,
byten	byte,
allmän	general,
river	tear,
avled	died,
någon	someone,anybody,
kriterier	criteria,
ses	be,
ser	sees,
förhöjd	enhanced,elevated,
sex	six,
sed	sed,
psykologiska	psychological,
uppkomsten	onset,
lyckas	successful,succeed,
järnväg	railway,rail,
sen	then,since,
något	any,something,
sorters	kinds,kinds of,
trey	trey,
guinea	guinea,
neutralitet	neutral,
fission	fission,
kejsarens	emperor,the emperor's,
stärkelse	starch,
alqaida	al-qaida,al-qaeda,
rita	draw,drawing,
europe	europe,
europa	europe,european,
påverkar	affecting,
giftermål	marrige,marriage,
medveten	aware,
avvikelser	abnormalities,deviations,derivations,
medvetet	consciously,conscious,
möts	meets,meet,
fame	fame,
stadsdel	district,
demografiska	demographic,demographical,
forskare	scientists,
bästa	the best,best,
medicinering	medication,
förändring	change,
bäste	best,
messias	messiah,
stå	stand,
kopia	copy,
samma	same,
transeuropeiska	transeuropean,
upprättades	was established,
krisen	crisis,the crisis,
kriser	crises,
church	church,
allierade	allied,allies,
decennium	decade,
sommaren	summer,
koalition	coalition,
mått	measurements,measurement,
väntade	waited,
tillväxt	growth,
kyrilliska	cyrillic,
upprättas	established,establish,
utsläpp	emission,emissions,
pågår	underway,
föranledde	brought about,led,
beskrevs	was described,described,
skönhet	beauty,
östafrika	east africa,
fire	fire,
taube	taube,
hovrätten	court of appeals,the court of appeal,
fritz	fritz,
uppleva	experience,
fritt	free,
föreningar	compounds,
systematik	systematic,
framträder	stand,appear,
projekt	project,
budget	budget,
feminism	feminism,
individerna	subjects,
bestående	comprising,lasting,
brottslighet	criminality,crime,
pressen	press,the pres,
föreställa	imagine,
arbete	work,
von	von,
owen	owen,
motors	motor,
teoretisk	theoretical,
erkänna	recognize,
slöts	signed,
lokaler	facilities,place,
korruptionsindex	corruption perceptions index,corruption index,
arbeta	working,
kritiker	critics,
barney	barney,
gärning	deed,
möjlighet	oppertunity,possibility,
omvandlas	converted,
omvandlar	converts,
skalet	shell,the shell,
barnen	children,
arméer	armies,
kritiken	criticism,the criticism,
laddning	charge,
kategoriavlidna	category deceased,
snarare	rather,
republiken	the republic of,the republic,
skapade	created,
debatten	the debate,
kring	on,around,
ledarskap	leadership,
fyra	four,
vargar	wolves,
euro	euro,
normala	normal,
krigsmakt	military power,armed forces,
person	person,
kelly	kelly,
johan	johan,
kontakter	contact,contacts,
finansiellt	financial,
sannolikhet	probability,
tunnelbana	subway,
stränder	beaches,
släppas	released,be released,
telegram	telegram,
stockholms	stockholm's,
finansiella	financial,
kontakten	connector,the contact,
mandat	mandate,
fascistiska	fascist,fascistic,
rebecca	rebecca,
festivalen	the festival,
symbolisk	nominal,symbolic,
nordväst	north west,
festivaler	festivals,
jönssonligan	jönssonligan,
tomas	tomas,
hennes	her,
format	format,shaped,
turnéer	tours,
teologiska	theological,
melker	melker,
avvisar	reject,
samarbete	co,
ivar	ivar,
västsahara	western sahara,
samarbeta	co,
da	da,
funnit	found,
skarp	sharp,crisp,
utlösa	trigger,
informationen	the information,
patrick	patrick,
ivan	ivan,
ulrich	ulrich,
lenin	lenin,
saknar	lacks,
saknas	missing,
användbar	useful,
utvecklades	developed,
avskaffade	abolished,absolished,
nåd	mercy,grace,
wallenstein	wallenstein,
öka	increasing,
brasilianska	brasilian,brazilian,
trafiken	the traffic,
turnerade	toured,
religion	religion,
riksförbundet	national association,
säger	said,says,
be	be,
norra	north,northern,
ugandas	uganda,
bl	bl,
vagnar	carts,carriges,
bo	living,
bk	bk,
plocka	pick,
engelska	english,
bokstav	character,letter,
ordning	system,
engelske	english,
by	by,village,
källor	source,
ideologin	ideology,the ideology,
bosättningar	settlements,
patrik	patrik,
soldaterna	soldiers,the soldiers,
dagligen	day,daily,
gemenskaperna	communities,community,
aggressiv	aggressive,
arméerna	armeerna,
stuart	stuart,
för	of,
papper	paper,
texterna	text,
inte	not,
inta	taken,
colorado	colorado,
syret	the oxygen,oxygen,
hemingway	hemingway,
efterföljande	subsequent,
spridas	spread,disseminated,
kraven	the demands,requirements,
popsångare	pop singer,
uppkallad	named,
orsaken	cause,
förlaget	publisher,
seger	victory,
veckor	weeks,
kategorimusikgrupper	category of music groups,
dröja	take,
utbröt	erupted,broke out,
samerna	sami,
knuten	tied to,knot,
fattigdom	poverty,
förbindelse	connection,
européerna	europeans,
poster	positions,post offices,
rörlighet	mobility,movement,
pastor	pastor,
begreppen	the concepts,terms,
begreppet	the term,concept,
posten	post,
atom	atom,
kritisk	critical,
line	line,
lovade	promised,
lina	lina,
dröm	dream,
fader	father,
cia	cia,
ut	out,
drogmissbruk	drug,
eddie	eddie,
ur	out,
konventionella	conventional,
distrikt	district,
uk	uk,
protestantiska	protestant,
lågt	low,
testamente	testament,will,
professor	professor,
översvämningar	flooding,
nämner	mentions,
pernilla	pernilla,
diverse	miscellaneous,
utbyggt	develpoed,built,
makedonska	macedonian,
nationalism	nationalism,
inblandning	incorporation,involvement,
iis	ii's,
händelsehorisonten	the event horizon,
räkna	count,
värld	world,
edwards	edwards,edward's,
são	sao,
skrivits	down,
innehåller	contains,
nordafrika	north africa,
innehållet	content,
matematiker	mathematician,
siffror	figures,numbers,
individuella	individual,
besegra	defeat,
dominerades	was dominated,dominated,
radikala	radical,
djurgårdens	djurgården's,
lucia	lucia,
ägnar	spend time,spends time,
konstantinopel	constantinople,
riskerar	risks,
springsteen	springsteen,
radikalt	radically,
slås	is hit,
alltså	therefore,really,
land	country,
passagerarna	passengers,the passengers,
uppträdande	performance,conduct,
symtom	symptoms,symptom,
age	do,age,
texten	text,the text,
sawyer	sawyer,
texter	texts,
majs	corn,
förväntas	expected,
persbrandt	persbrandt,
släpptes	released,was released,
alltför	all too,way too,
bakåt	backwards,reverse,
turkisk	turkish,
dyraste	most expensive,
hamnar	lands,ports,
young	small,
listade	listed,
dickinson	dickinson,
dancehall	dancehall,
sent	late,
garden	garden,
märken	sign,
kedjan	chain,the chain,
palestinier	palestinians,
kommunistiska	communistic,communist,
flöde	feed,
drogen	the drug,drug,
känner	knows,
överleva	survival,
tillhörande	associated,belonging to,
magic	magic,
påverka	impact,influence,
harbor	harbor,
eva	eva,
tre	three,
jobbet	work,the job,
romerska	roman,
överlevt	survived,
romerske	roman,
opinionen	opinion,
innebörden	meaning,the significance,
leonardo	leonardo,
bolsjevikerna	bolsheviks,the bolsheviks,
natur	nature,
regelbundna	regular,
ställde	set,
förhållandevis	relatively,
legitimitet	legitimacy,
victor	victor,
antog	adopted,
index	index,
expressen	expressen,
anton	anton,
praktiken	effectively,
indiens	indias,
suveräna	terrific,
möjliggör	enables,enable,
birk	brik,birk,
indian	indian,
ledande	conductive,leading,
stadskärna	town,
led	suffered,step,
lee	lee,
lyckades	managed,succeeded,
upphovsrätten	copyright,
sålunda	thus,
leo	leo,
lev	lev,
hälsa	health,
talang	talent,
begravd	buried,
motorvägarna	highways,the highways,
solen	sol,
tegel	brick,
casino	casino,
titanic	titanic,
förutsätter	assume,requires,assumes,
tillkom	hold back,resided,
insulin	insulin,
högsta	highest,
opinion	opinion,
artisterna	artists,
huvudvärk	headache,
emot	vis,
förlora	lose,
oxenstierna	the oxenstierna,oxenstierna,
mening	sentence,
indianerna	the indians,indians,
anatolien	anatolia,
andreas	andreas,
varmare	warmer,
rico	rico,
illegal	illicit,
hemlig	secret,
elever	students,
godkänna	approve,
klaviatur	keyboard,
orkester	orchestra,
projektet	project,
existerade	existed,
författning	constitution,
samspel	teamwork,
ytterst	highly,
överlevande	survivors,
villor	villas,
indianska	native american,
lokalt	locally,local,
bidraget	grant,
advokat	bar,
ortodoxa	orthodox,
lokala	local,
peka	point,
sekel	centuries,
upprätthålla	maintaining,
process	process,
klassisk	classical,
etta	number one,first,one,
syre	oxygen,
high	high,
tryckta	printed,
hercegovina	herzegovina,
sydöstra	south east,
halmstad	halmstad,
frågor	questions,
saknade	missed,missing,
delad	divided,
övergrepp	assault,abuse,
latinska	latin,
hormoner	hormones,
delas	shared,divided,
delar	proportions,parts,
delat	shared,
sydvästra	southwest,southwestern,
kriminella	criminal,
amerika	american,america,
djurens	the animals,
profeten	prophet,the prophet,
insatser	action,
regeringsmakten	government power,
väckt	brought,awaken,
slutsatser	conclusions,
spelen	the games,
lundgren	lundgren,
nancy	nancy,
napoleons	napoleon's,napoleon,
byggnadsverk	building,
borde	should,
handboll	handball,
diskar	disks,
möjligt	possible,
hårdast	hardest,the hardest,
universiteten	universities,the universities,
frånvaro	absent,absence,
hunnit	had time to,
universitetet	the university,university,
solvinden	the solar wind,solar wind,
västerbottens	västerbottens,west bothnia,
eliten	the elite,elite,
uppdelat	split,
tecknet	the sign,sign,
uppdelad	divided,split,
puerto	puerto,
beståndsdelar	constituents,elements,
ovanlig	rare,uncommon,
bekant	known,acquaintance,
bryter	breaks,
hemmaplan	home,
dock	nevertheless,however,
utgår	deleted,
rotation	rotation,
huvuddelen	bulk,
sönder	broken,
peking	beijing,peking,
välfärd	wealth,welfare,
intressen	interests,
fortsätta	remain,continue,
smallwood	smallwood,
fördrevs	was banished,
överföras	transfer,transferred,
books	books,
intresset	the interest,
frac	fraction,
banan	banana,
etymologi	etymology,
matrix	matrix,
borderline	borderline,
trycktes	was published,printed,
enskilda	individual,
anledningen	therefore,
umgänge	intercourse,
kapitalismens	capitalism,capitalism's,
marxistiska	marxist,
bekräftades	was confirmed,
fram	out,
undertecknades	signed,
redskap	device,tool,
egenskaperna	the qualities,properties,
statschef	head of state,
påverkats	affected,
melankoli	melancholy,
uppe	up,
förts	brought,
tempererat	temperate,
dubbel	double,
liggande	placed,
kompositör	composer,
krävt	required,
våldsam	violent,
krävs	needs,requires,
david	david,
blanda	mix,
profeter	prophets,
krets	sphere,circuit,
helst	rather,anyone,
hussein	hussein,
kräva	require,
skillnad	difference,unlike,
playstation	playstation,
åring	year old,years,
komplicerade	complex,
jesus	jesus,
användningsområden	possible use,applications,
schweiziska	swiss,
muhammad	muhammad,
nordkoreanska	north korean,
studerade	studied,
värdefulla	valueable,value,
artiklar	items,
festival	festival,
system	system,
bygget	construction,
syster	sister,
hebreiska	hebrew,
tränga	permeate,cut in,
teatern	the theater,
blivit	become,was,
utbyggnad	development,expansion,
havet	sea,
pristagare	laureate,
utländska	foreign,
haven	the seas,
visdom	wisdom,
hampa	hemp,
samverkar	co,
roberto	roberto,
stewie	stewie,
roberts	roberts,
reagans	reagan's,reagan,
troende	believers,faithful,
samverkan	co,
jonatan	jonatan,
räcker	enough,sufficient,
användaren	the user,user,
producent	producer,
förslag	proposed,
flygplats	airport,
element	elements,
kritiskt	critical,
instruktioner	instructions,
mills	mills,
filosofin	philosophy,the philosophy,
sinatra	sinatra,
kritiska	critical,
best	best,
linda	linda,
viss	certain,some,
finsk	finnish,
slutsatsen	concluded,the conclusion,
säkert	securely,
nät	web,
trosbekännelsen	creed,
detta	that,
vardagen	the weekday,everyday life,
kvinnliga	female,
visa	see,
uppror	rebellion,
flyga	fly,
förutsättningarna	prerequisites,conditions,
medan	while,
framgår	will be seen,is shown,
synliga	visible,
våren	spring,the spring,
bokstaven	the letter,character,
face	face,
synligt	seen,
befolkningens	population,
närmade	approached,
brev	letter,
beteende	behaviour,
uppdelade	divided,
manchester	manchester,
tyvärr	unfortunately,
hopp	hopes,hope,
fursten	prince,
östfronten	eastern front,the east front,
samisk	sami,
jan	jan,
religionens	religion,religion's,
liksom	and,
jah	jah,
jag	i,
skarsgård	cut farm,skarsgård,
ilska	anger,
abba	abba,
parlamentet	the parlament,parliament,
lägger	put,lies,
fotbollsspelare	football player,footballers,
lucky	lucky,
generalen	the general,general,
bonde	farmer,
parlamenten	parliaments,
meter	meters,meter,
tidigaste	earliest,
britterna	the brits,british,
h	h,
rowling	rowling,
effekterna	the effects,effects,
iranska	iranian,
rymmer	holds,
guvernör	governor,
myndigheterna	the authorities,the authoroties,
debuterade	debut,debuted,
michail	michail,
priser	rates,prizes,
avlidit	died,
priset	the prize,rate,
kronisk	chronic,
uppträdde	perform,occurred,
lämplig	suitable,
freddy	freddy,
sköt	shot,
vietnams	vietnam's,vietnam,
författarskap	the writer,authorship,
sjöng	sang,
upprättandet	establishment,establishing,
längst	at,farthest,longest,
sjönk	sunk,sank,decreased,
balansen	balance,the balance,
varning	warning,
kategorisvenskar	category swedes,
striden	battle,
finalen	final,
bolivias	bolivia,bolivia's,
strider	battles,
bilar	car,cars,
ende	only,
förklaringar	explanations,
kedjor	chains,
islamiska	islamic,
ett	a,
marknaden	the market,market,
figuren	the character,figure,
beläget	located,base,
fåglar	birds,
egypten	egypt,
norge	norway,
etc	etc.,
marknader	markets,
ogillade	disliked,
belägen	disposed,
utövade	exerted,exercised,
tätbefolkade	densely populated,populated,
ekvatorn	equator,the equator,
religiösa	religious,
botten	bottom,
co	co,
dör	dies,
ca	cirka,approximately,
mengele	mengele,
cd	cd,
stabila	stable,
cp	cp,
öst	east,
dök	appeared,dove,turned,
antal	number,
jussi	jussi,
keltiska	celtic,
företaget	the company,
moraliskt	morally,moral,
överallt	in all,everywhere,
kombination	combination,
växt	plant,
genetik	genetics,
moraliska	moral,
företagen	the companies,
antas	assumed,
antar	adopting,
regelbundet	regularly,
molekyler	molecules,
tvungna	forced,forced to,
undervisningen	teaching,the education,
sänts	sent,
atlanta	atlanta,
haile	haile,
mandatperiod	term of office,
långsamma	slow,
tjorven	tjorven,
rikets	its,the realms,
demokrati	democracy,
aktivitet	activity,
vd	ceo,
ondskan	the evil,
förlopp	process,developments,
omnämns	mentioned,is mentioned,
vi	we,
ryssland	russia,
vm	world championship,vm,
lust	loss,
vs	vs,
flickor	girls,
skapare	creator,
föreligger	exist,
sitt	its,
slovenska	slovenian,
spela	play,
tupac	tupac,
armé	poor,
känt	known,
juan	juan,
medeltida	medival,medieval,
foundationthe	the foundation,
huden	skin,
romance	romance,
känd	known,unknown,famous,
terrorism	terrorism,
flesta	most,
ball	ball,
columbia	columbia,colombia,
sade	said,
framförde	performed,presented,
anordnas	provided,arranged,
anfield	anfield,
ikea	ikea,
sjukhus	hospitals,
diabetes	diabetes,
representera	represents,represent,
mänskligt	human,
klubbarna	the clubs,
väger	weighs,weight,
vägen	the road,
ledde	resulted,
ledda	led,
uno	uno,
versaillesfreden	versailles peace,treaty of versailles,
vägarna	paths,
gatan	the street,
paus	pause,paus,
aktuell	current,
renässansen	the renaissance,renaissance,
paul	paul,
pappa	dad,
installera	installing,
förknippas	associated to,
planeter	planets,
frågan	issue,the question,
englands	england's,
planeten	planet,the planet,
kosovos	kosovo,
filmens	the film's,
framtid	future,
förknippad	associated,
motorvägen	highway,
government	government,
ledarna	the leaders,conductors,
gul	yellow,
dess	its,
arbetarklassen	working class,the working class,
tillverkning	production,
pressas	pressed,
följeslagare	companions,companion,
lät	had,
emma	emaa,emma,
lär	teach,learn,
aktiebolag	stock company,
vallhund	herding dog,
stadsbild	cityscape,
amazonas	the amazon rainforest,amazon,
symptomen	the symptoms,
högskolan	hogs school,university,
flotta	fleet,
län	state,
tackade	thanked,said/thanked,
bredare	broad,
miniatyr|	miniature,
filmografi	filmography,
anarkismen	the anarkism,anarchism,
trotskij	trotskij,trotsky,
lägsta	lowest,
stannar	stays,
transport	carriage,transportation,
skriftliga	written,
ockupation	occupation,
februari	february,februari,
behandlades	treated,
flitigt	actively,frequent,
tänkandet	thinking,the way of thinking,
dags	time,
naturlig	natural,
kollektivtrafik	public transport,
ateist	atheist,
svaga	weak,
förklaringen	the explanation,statement,
biologi	biology,
överlevnad	survival,
östberlin	east berlin,
svagt	weak,
gandalf	gandalf,
smärta	pain,
vargen	the wolf,
användande	use,
kontinenten	the continent,
må	mon,
erövrade	conquered,
höger	right,
blodiga	blooded,bloody,
angeles	angeles,
kontinenter	continents,
warner	warner,
solsystemets	solar system,
hittills	date,
släpper	release,releases,
upplösningen	dissolution,disbandment,
sekelskiftet	turn,
planetens	the planets,
kristus	christ,
lund	grove,
mera	more,
ting	matters,
peters	peters,
skola	school,
fläckar	stain,
bedöms	expected,
överbefälhavare	commander-in-chief,supreme commander,
tina	defrost,thaw,
radioaktiva	radioactive,
samlingar	collection,
förre	pre,
uppvisade	showed,
apollo	apollo,
radioaktivt	radioactive,
svält	starvation,starvations,
återkommer	will return,
society	society,
volvo	volvo,
ruset	the fuddle,intoxication,
stormakt	great power,
monument	monument,monuments,
inrättades	established,were implemented,
distribution	distribution,
distriktet	district,
leukemi	leukemia,
heter	units,
guy	guy,
utnyttjar	using,
utnyttjas	utilized,used,
skilsmässa	divorce,
separerade	separated,
broder	brother,
vitryssland	belarus,
månader	months,
sharia	sharia,
öga	eye,
distinkta	distinct,
särskilt	in particular,especially,
relationen	the relation,ratio,
månaden	the month,months,
modernistiska	modernistic,modernist,
bröd	bread,
övergång	transition,
francisco	fransisco,
uttalade	spoke,
tider	times,
förhandlingar	negotiations,
bröt	broke,
tiden	time,
inspiration	inspiration,
syskon	siblings,
mozart	mozart,
sänker	lowers,lower,sinks,
tredje	third,
jordbävning	earthquake,
provinser	provinces,
kommersiell	commercial,
nederländska	netherlands,dutch,
brevet	the letter,letter,
näsan	the nose,nose,
child	child,
elisabeth	elisabeth,
bosniska	bosnian,
tätort	urban,conurbation,
invadera	invade,
preussen	prussia,
konsekvenserna	impact,
smålands	småland,
bäst	best,
atlanten	the atlantic ocean,
bibel	insulin,bilble,
spel	game,
edward	edward,
nervsystemet	nervous system,the nervous system,
nödvändigt	neccessary,necessary,
ale	ale,
mördade	murdered,
konsekvent	consistent,consistency,
grönsaker	vegetables,
golvet	the floor,floor,
främste	chief,premier,
geologi	geology,
jacob	jacob,
skolor	schools,
innefattar	comprises,includes,
uttryck	expression,
upphörde	ceased,
estland	estland,estonia,
jamaica	jamaica,
ständerna	the cities,
galax	galaxy,
horn	horns,horn,
colorblack	color black,
alltsedan	since,
förbättringar	improvement,
eurovision	eurovision,
bakgrunden	background,
vidsträckta	broad,
kraftfull	forceful,
tolv	twelve,
bidrag	contribution,contributions,
vampyr	vampire,
cyklar	bicycles,cycles,
bidrar	contributes,
petra	petra,
musikalen	the musical,
räddar	saves,rescues,
bortgång	passing,death,
pluto	pluto,
rapporterar	reports,
norstedt	norstedt,
begått	committed,
olsson	olsson,
studeras	studied,is studied,
studerat	studied,
interstellära	interstellar,
regerande	ruling,
hänvisade	referred,
förblir	remains,
stoft	dust,
träda	esterified,emerge,fallow,
placerades	placed,
akc	akc,
underverk	wonders,
diameter	diameter,
järnmalm	iron ore,
fastställdes	confirmed,set,
bro	bridge,
läkemedelsverket	food and drug administration,
faktiska	actual,
total	total,
bra	good,
stått	stood,
sarah	sarah,
ätten	the dynasty,dynasty,
negativa	negative,
foster	fetal,
indiana	indiana,
negativt	negative,
supportrar	supporters,
ifall	if,
förebyggande	preventive,
giovanni	giovanni,
award	award,
riksväg	national highway,
nku	nku,
alces	alces,
lissabonfördraget	treaty of lisbon,lisbon treaty,
kurderna	kurds,
absorberas	absorbed,
friheten	freedom,liberty,
beväpnade	armed,
fascismen	the fascism,fascism,
dokument	documents,
era	yours,era,
transparency	transparency,
specialiserade	specialized,special,
klorofyll	chlorophyll,cholophyll,
vietnamesiska	vietnamese,
gloria	gloria,
vackra	beautiful,fine,
felaktiga	false,
ekonomiskt	economically,economical,
sommar	summer,
indien	india,
indier	indians,
enhet	unit,entity,
valborg	may day,valborg,
utlandet	abroad,
gotlands	gotland's,gotland,
ansluter	connects,
firas	celebrated,celebrate,
firar	celebrates,celebrate,
gillar	like,likes,
halland	halland,
beach	beach,
sammansatt	composed,compound,
biografer	movie theaters,
kategorieuropas	category europe,
lag	law,act,
koreakriget	korean war,the korean war,
visste	did,
tjäna	profit,
biografen	movie theater,cinema,
law	law,
orden	the words,words,
medlemsstat	member state,
vänsterpartiet	leftist party,left wing party,
lämningar	remnants,
green	green,
massmedia	media,
livets	life,life's,
ordet	word,
order	order,
arbetslöshet	unemployment,unemplyment,
natten	overnight,
office	office,
sovjet	soviet,
diagnos	diagnostics,
exempel	example,
ramadan	ramadan,
söderut	south,
blandning	mix,mixture,
japan	japan,
bidra	contribute,
straff	punishments,
lagets	substrate,the team's,
fragment	fragments,
vanligtvis	usually,generally,
ämne	substance,
band	band,
fredsbevarande	peace,peacekeeping,
bana	course,web,
they	they,
spelningen	the gig,
bank	bank,
ansvariga	charge,
huvudartikel	main article,
helvetet	hell,
dåliga	poor,bad,
diskuteras	discussed,
knutpunkt	hub,
dåligt	poor,
område	area,
carlos	carlos,
erbjöd	offered,
germanska	germanic,germanian,
inflytandet	the influence,influence,
koldioxid	carbon dioxide,
däggdjur	mammalian,
rummet	room,
kejserliga	imperially,imperial,
asteroidbältet	asteroid belt,the asteroid belt,
daniel	daniel,
levnadsstandarden	the standard of living,standard of living,
trafik	traffic,
bruttonationalprodukt	gross national product,bnp,
oskar	oskar,
vete	wheat,
klimatet	climate,
veta	out,
sedermera	subsequently,since,
veto	veto,
standard	standard,
tillbaka	back,
berör	affecting,affect,concerns,
amadeus	amadeus,
ange	set,
sprit	alcohol,
väldiga	immense,mighty,vast,
förefaller	appears,
professionell	professional,
väldigt	very,
förmågan	the ability,
personerna	subjects,
funktioner	features,
önskar	desired,wish,
önskan	desired,
another	another,
statskupp	coup,
ingmar	ingmar,
drabbade	affected,
begränsas	limited,
begränsar	limit,limits,
ingen	no,
begränsat	limited,restricted,
sång	song,
lidande	sufferer,
växthusgaser	greenhouse gas,
inget	not,no,
john	john,
begränsad	restricted,
medborgare	citizens,
antisemitismen	anti-semitism,
äter	eat,eats,
varifrån	from which,
albert	albert,
åland	Åland,
kvarvarande	remaining,
persson	persson,
bojkott	boycott,
kraftverk	power plant,
trupp	troops,troop,
finska	finnish,
militära	military,
nedan	below,
symboliserar	symbolizes,
binda	bond,
sonen	the son,
scener	scenes,
används	use,
scenen	stage,
binds	bind,
iron	iron,
byggts	built,
minut	minute,
använde	used,
använda	using,
årens	the year's,years,
skolorna	schools,the schools,
mannen	art,the man,
noterade	note,
onani	masturbation,
fåglarna	birds,
omvandling	transformation,
framtida	future,
koloniala	colonial,
småningom	eventually,
kalendern	calendar,calender,
stavning	spelling,
magnus	magnus,
höjd	height,
sjukvård	healthcare,
aftonbladet	aftonbladet,newsweek,
lades	put,
anatomi	anatomy,
närvaro	attendance,presence,
verkat	worked,seemed,
verkar	acting,seems,
maiden	maiden,
bruce	bruce,
utställning	display,exhibition,
skansen	forecastle,
fjädrar	feathers,
verkan	effect,
flygplatsen	airport,the airport,
aminosyra	amino acid,
vägg	wall,
eviga	eternal,
ägda	owned,
freja	joe,
ägde	was,owned,
bortom	beyond,beyond the,
läran	the teaching,
evigt	forever,
misslyckade	failed,
förväxla	confuse,mistake,
effekten	the effect,effect,
mitten	middle,
damer	ladies,
lewis	lewis,
hinduiska	hindu,
vanligen	usually,typically,
tilläts	was allowed,
effekter	effects,
fortplantning	reproduction,
vätet	hydrogen,the hydrogen,
sättet	manner,the way,
 kilometer	kilometer,
sätter	place,puts,
estetiska	aesthetic,
ambassad	embassy,
kejsar	emperor,
inställning	attitude,setting,
målvakt	goalee,goalkeeper,
kontinuerlig	continuous,
imperium	empire,
dj	dj,
di	di,
de	the,they,
dc	d.c.,
sverigedemokraterna	sweden democrats,
stalins	stalins,
watson	watson,
människorna	men,
orolig	worried,
riktningen	direction,denomination,
du	to,you,
dr	doctor,
sattes	was added,
peyton	peyton,
offret	the victim,
runt	around,
spridningen	proliferation,the spread,
konst	art,srt,
sentida	recent,
splittrades	split,
offren	victims,
tyngre	heavy,heavier,
fågelarter	species of bird,
viktigt	important,
libanon	lebanon,
kurdiska	kurdish,
vanlig	ordinary,normal,
utförd	completed,performed,
utföra	perform,out,
förena	combine,unite,combining,
väsen	being,
historiens	historys,
präglats	been characterized,
utfört	done,
massiva	solid,
utförs	out,
sexuell	sexual,
djuret	the animal,animal,
fornnordiska	ancient nordic,old norse,
månarna	moons,
fångenskap	captivity,
piratpartiet	pirate party,
djuren	animals,
materialet	the material,material,
smaken	the flavour,flavor,
osmanska	osmanian,
komplikationer	complications,
we	we,
självständigheten	independence,
förkortningar	abbreviations,
miljö	environment,
jämförelse	comparative,comparison,
huvudsakligen	generally,primarily,
militären	military,the military,
garanterar	ensures,guarantees,
kännetecknas	is characterized,
cox	cox,
startade	started,
kommer	is,
brad	brad,
målningen	milling,the painting,
vecka	week,
graviditeten	the pregnancy,
kännetecken	distinction,sign,
thierry	thierry,
fångar	captures,prisoners,
chrusjtjov	khrushchev,chrusjtjov,
genomför	implement,out,
tony	tony,
slaveriet	slavery,
smith	smith,
japans	japans,
patienten	patient,the patient,
tids	time,
lösning	solution,
framträdande	apperance,
hitlers	hitlers,
patienter	patients,
klubblag	club team,
attacken	the attack,attack,
attacker	assaults,
fest	party,fest,
juridik	law,
drottningen	queen,the queen,
frekvens	frequency,
förstnämnda	first named,
bulgariens	bulgaria,
fromstart	starting from,
vagn	carrige,
johansson	johansson,
påstådda	alleged,
kupp	kupp,coup,
aik	aik,
anhängare	supporters,
nordöstra	nordeastern,northeast,
spanjorerna	spaniards,the spaniards,
gärdestad	nugent,
have	have,
moldavien	moldova,
deltagarna	the participants,participants,
jordbruk	agricultural,
påverkades	was affected by,affected,
själva	self,actual,
våg	road,wave,
patent	patent,
datorer	pc,
bergskedjor	mountain ranges,
från	from,
självt	itself,
utgivna	published,
bunny	bunny,
andelen	the share,the proportion,
producerades	produced,
raid	raid,
hann	did,reached,
saddam	saddam,
balkan	the balkans,
sexualitet	sexuality,
delstater	states,
delstaten	the state,
nervosa	nervosa,
hans	his,
bilen	the car,car,
koncentrerad	concentrated,
aspekter	aspects,
rörelsen	movement,
rör	touches,
styrkorna	forces,
mamma	mother,
monaco	monaco,
rörelser	movement,
röd	red,
thc	thc,
skottland	scotland,
gärningsmannen	culprit,
newton	newton,
kall	cold,
nästan	almost,close,
kroppens	the body's,the bodies,
goda	good,
enades	agreed,
kalender	calendar,calender,
upptäckte	discovered,
swahili	swahili,swahilli,
så	as,so,
distributioner	distributions,
snus	snuff,
havets	the seas,sea,
skick	state,condition,
kvinnan	female,
samfund	communities,order,
plasma	plasma,
född	born,
maya	maya,
föda	feed,
återgick	returned,returning,
skadorna	damages,damage,
arab	arab,
fusion	fusion,
indianer	indians,
föds	born,
everton	everton,
picasso	picasso,
hepatit	heptatitis,
acceptera	acceptable,
årlig	yearly,
indelning	the subdivision,classification,
indelningen	division,subdivision,
dahlén	dahlén,
xbox	xbox,
gandhi	gandhi,
transkription	transcript,
sixx	sixx,
avsätta	depositing,
bort	away,
born	born,
presidentvalet	presidential elections,presidential election,
borg	tower,castle,
bord	table,
kungar	kings,
humor	humor,humour,
territorierna	territories,
purple	purple,
serbiens	serbias,
siffran	number,figure,
columbus	columbus,
stadsdelarna	districts,
vägar	roads,
bevara	preserve,preserving,
post	week,
slovakien	slovakia,
vunnit	won,
banker	banks,
olika	different,variety,
jacques	jacques,
återfinns	found,is rediscovered,
samer	sami,
karlsson	karlsson,
epicentrum	epicentre,epicenter,
fängslade	inprisoned,imprisoned,
blivande	prospective,future,
effekt	effect,power,
gemenskapen	the collective,community,
way	way,väg,
was	was,
war	war,
expansionen	expansion,the expansion,
hypotes	hypothesis,
skiljas	separated,separate,
motorvägar	highways,
inträffar	occur,
inträffat	occurred,
partiledare	party leader,
emil	emil,
reser	travels,
studierna	the studies,
mtv	mtv,
finansiering	financing,
litterär	literary,
långvarig	long,
träning	training,
erövra	conquer,
engagerade	dedicated,engaged,
moore	moore,
utomlands	abroad,
tesla	tesla,
xiis	xii,
efter	after,
bilderna	the pictures,
moln	cloudy,
empati	empathy,
toppen	the top,
cellerna	cells,the cells,
möta	meet,face,
förmåga	abilities,ability,
janukovytj	janukovytj,yanukovych,
möte	meeting,
arkitekter	architects,
test	test,
götaland	götaland,
konservatism	conservatism,
mött	met,
femton	fifteen,
tottenham	tottenham,
räknat	calculated,counted,
reglerar	regulates,controls,
regleras	is regulated,controlled,
rätter	dishes,
omgivande	surrounding,surounding,
rätten	right,the court,
solens	solar,
bergmans	bergman's,bergmans,
dance	dance,
uppfanns	was invented,invented,
global	global,
datum	date,
redaktör	editor,
osäker	unsure,
lider	suffering,suffers,
utkämpades	fought,
förhistorisk	prehistorian,
afrikaner	africans,
heller	nor,
rådet	council,
igelkott	hedgehog,
zone	zone,
vattenånga	steam,water vapour,
vänder	turn,face,
division	division,
hannah	hannah,
uttrycka	express,
lättare	light,easier,
hannar	males,
uttryckt	expressed,
enskilt	individually,single,
salvador	salvador,
stycken	pieces,
gud	god,
konstnärlig	art,artistic,
sätt	manner,way,
hisingen	hisingen,
levnadsstandard	standard of living,
frigörs	released,is released,
ljuset	the light,light,
säte	seat,
formella	formal,
litterära	literary,literal,
templet	temple,
revolution	revolution,
alfa	alpha,
cosa	cosa,
engagerad	dedicated,engaged,
invandrade	immigrated,immigrant,
sköttes	operated,handled,
mål	case,
motsatte	opposed,
midsommar	midsummer,
stimulera	stimulate,stimulating,
motsatta	opposite,
yorks	yorks,
ungdomar	youths,
tidig	early,
ingick	were included,was,
kosmiska	the cosmic,cosmic,
uniform	uniform,
fastigheter	real estates,properties,
utspelar	takes place,set,
versionen	edition,the version,
gener	genes,
oerhörd	tremendous,
marxismen	marxism,
kärlek	love,
påstås	claimed,
påstår	states,claims,asserts,
genen	the gene,
oerhört	tremendously,
tillträde	access,
antarktiska	antarctic,
sistnämnda	later,last,
kemi	chemistry,
franklin	franklin,
ponny	pony,
vinnare	win,winner,
ekr	ekr,ad,
marken	soil,
vapnet	the weapon,
spridit	spread,disseminated,
ukrainas	ukrainian,
vapnen	weapons,the weapons,
förteckning	listing,
kärnkraftverk	nuclear power plant,
presenterar	presents,present,
upprättade	established,prepared,
äktenskapet	marriage,
super	super,
stabilitet	stability,
live	live,
regel	rule,
territoriet	territory,
angels	angels,
överhuvudtaget	in general,
fransmännen	the french,
parallellt	parallel,
rivalitet	rivalry,
snabbt	fast,quickly,
enda	only,
målvakten	the goalkeeper,
zarathustra	zarathustra,
ämnena	subjects,the elements,
närmar	close,closing,close in,
varför	therefore,why,
norrköpings	norrköpings,
feministiska	feminist,
snabba	rapid,
löner	salaries,
ibm	ibm,
ibn	ibn,
interaktion	the interaction,interaction,
frukt	fruit,fruits,
can	cancer,
erbjuder	offers,
heart	heart,
några	few,a few,
december	december,
nobels	nobel's,
influensavirus	flu virus,influenza,
gentemot	towards,against,
abort	abortion,
uppstår	occur,
genomgått	experienced,passed,
kritiserar	criticize,
ligan	league,
pojke	boy,
uppskattades	was appreciated,
betydelse	importance,significance,
kopplingar	connections,
perserna	the persians,
southern	southern,
framgångarna	successes,
göteborgs	gothenburg,gothenburgs,
gräns	border,
ungern	hungary,hungaria,
förutsättning	provided,prerequisite,
romarna	romans,the romans,
flyttas	moved,
flyttar	move,
kurt	kurt,
kurs	course,
ukrainska	ukrainian,
rekordet	record,the record,
maktens	the powers,forces,the power's,
landshövding	county governor,
ingripa	act,
ganska	quite,
ättlingar	descendants,
magnetfält	magnetic,magnetic field,
generalguvernören	general governor,
linnés	linnaeus,
fält	field,
skabb	mites,scabies,
levde	lived,survived,
utnämndes	was declared,appointed,
därifrån	from there,
bergskedjan	mountain range,the mountain group,
yngre	younger,
hals	throat,
varav	of which,
arton	eighteen,
varar	duration,lasts,
nog	enough,
författarna	the authors,writers,
förvaras	stored,is stored,
komponenter	components,
begränsa	limit,
not	note,
nou	nou,
rakt	straight,
now	now,
dödsstraffet	death penalty,
uppgörelse	settlement,agreement,
frihet	freedom,
språk	language,
främmande	undesirable,foreign,
antyder	indicates,
stockholm	stockholm,
januari	january,
drog	draw,pulled,drug,
aspergers	aspergers,
em	em,european championship,
el	el,
en	a,
citat	quote,
ej	not,
ed	ed,
utbrett	wide,widespread,
strålningen	radiation,
kroatiska	croatian,
et	et,
resultera	result,
fuglesang	fuglesang,
ep	ep,
premiärministern	prime minister,
er	you,
album	album,
teorier	theories,
återkommande	recurring,
videon	video,
hustrun	his wife,
kortare	shorter,
stallone	stallone,
punkt	item,point,
skära	carve,
välkänd	well-known,well known,
marina	marine,
betraktades	regarded,
åt	to,
böhmen	bohemia,
british	british,
domen	judgment,
allmänheten	public,general public,
arbetsgivare	employers,
blind	bank,blank,
xi	xi,
förändrats	changed,
derivatan	derivative,the derivative,
någorlunda	fairly,somewhat,
ring	ring,
xv	xv,
bergqvist	bergqvist,
våglängder	wavelength,
omtvistat	disputed,
konungarike	kingdom,
desmond	desmond,
sheen	sheen,
dessutom	moreover,furthermore,
satsningar	ventures,investments,
färre	less,
spelningar	gigs,
fascisterna	fascists,
delats	divided,been awarded,
television	television,
europeisk	european,
sidorna	the pages,pages,
utbyggda	expanded,
ändrades	changed,
kloster	monastery,
grundad	founded,based,
craig	craig,
statsminister	prime minister,
kairo	cairo,
grundat	founded,
utifrån	from,
grundar	bases,
grundas	is based,
anger	indicates,gives,
anges	is put at,specified,
befolkningstillväxt	population growth,
hjälp	using,help,
hör	include,hears,
form	form,
fortsatte	continued,
fortsatta	continued,
etiopiska	ethiopian,etiopian,
bönor	beans,
hög	high,
online	online,
skäl	reasons,
åtta	eight,
kategoriorter	category visited,
numera	now,
santiago	santiago,
successivt	successively,
bön	prayer,
bekostnad	detriment,expense,
dvärgar	dwarves,dwarfs,
glödlampor	light bulbs,
america	america,
på	on,
michelle	michelle,
lyfter	lift,lifts,
norrmän	norwegians,
nordligaste	northern,northernmost,
parlamentets	parliament,
runda	round,
orsaka	cause,
abraham	abraham,
skapats	was created,generated,
doktor	doctor,
kyrkorna	churches,the churches,
behåller	retain,
marocko	morocco,marocco,
colombo	colombo,
teori	theory,
perfekt	perfect,
mannens	man,
byggda	constructed,
rötter	roots,
varmblod	warmblood,
raúl	raul,
himmel	heaven,
huskvarna	huskvarna,
byggde	was,
dagbok	log,
sierra	sierra,
sydligaste	southernmost,most southern,
uppståndelse	resurrection,
helgdagar	holidays,
riddare	knight,
samuel	samuel,
gudarnas	the gods',gods,
ambitioner	ambitions,
folkomröstning	referendum,
marxistisk	marxist,
tävla	compete,
handlingar	actions,
drabbas	affected,
facupen	fa cup,fa-cup,
tvingade	forcing,
bushadministrationen	the bush administration,
länge	long,
storstäder	metropolises,cities,
tillfällig	temporarily,
osbourne	osbourne,
övergången	transition,
sport	athletics,sport,
katastrofer	disasters,catastrophes,
depressionen	the depression,depression,
konstaterade	established,
ladin	ladin,
depressioner	recessions,depression,
israels	israeli,israel's,
import	import,
kommunismens	communism,the communisms,
katastrofen	catastrophy,the catastrophy,
yta	surface,
ronja	ronja,
personlighet	character,personality,
flygande	flying,
männen	men,
utgivningen	the publication,the release,
verket	board,
rike	kingdom,
verken	plants,
utgavs	was published,published,
comeback	comeback,
samtal	conersation,call,
warhol	warhol,
representativ	representative,
bördiga	fertile,
placerad	disposed,
handlar	is,concerns,
kristinas	kristina's,crisis thawed,
propaganda	propaganda,
feminismen	feminism,
undersökning	study,
nils	nils,
placerar	places,
placeras	placed,
utnyttja	use,
avskaffande	elimination,abolition,
dömande	sentencing,judging,
regeringens	government,
lägenhet	apartment,appartment,
bomull	cotton,
östtyska	east german,
överlever	survives,
handlande	action,
långfilm	feature film,
oliver	olives,
välstånd	prosperity,
wien	vienna,
sker	is,
oden	node,oden,
knappt	barely,
socialdemokrater	social democrats,
dräkt	costume,outfit,
observera	note,observe,
utförda	formed,performed,made,
utförde	did,
elvis	elvis,
funnits	found,been,
konservativa	conservative,
ytan	the area,surface,area,
uefacupen	the uefa champions league,
rapporter	reports,
prinsessan	the princess,princess,
rapporten	report,
polens	polands,pole,
ordningen	the order,order,procedure,
ansikte	face,
tjeckien	czech republic,the czech republic,
eran	era,
tycker	thinks,
bevis	certificate,evidence,
finanskrisen	financial crisis,the financial crisis,
tänkande	thinking,
behandlade	treated,
kvarter	quarter,block,neighborhoods,
kenya	kenya,
västerländska	western,
katalanska	catalan,
helium	helium,
grundade	based,
infödda	natives,native,
slaget	the strike,type,
långt	long,
orsakade	caused,causing,
programvara	software,
media	media,
långa	long,
talmannen	president,
homosexualitet	homosexuality,
kromosom	chromosome,
pesten	the plague,plague,
lite	little,a little,
demens	dementia,
figurer	figures,
speciella	special,
offensiven	offensive,
begär	requests,request,
skivbolaget	record label,the record company,
acdc	ac/dc,
omfattande	large,
omfattar	include,
omfattas	comprise,subject,
speciellt	particularly,
omgående	immediately,immediate,
ekonomisk	economic,
tradition	tradition,
fredspris	peace prize,
skånes	scania,
erkänd	acknowledged,recognized,
flaggor	flags,
mynning	outfall,mouth,
forskarna	the scientists,
skandinaviska	scandinavic,
tydlig	clear,
framgången	success,the success,
samiska	sami,
eleverna	the pupils,the students,
lagerkvist	lagerkvist,
nazismen	nazism,
euron	the euro,euro,
malcolm	malcolm,
lade	laid,added,
ditt	your,
strävar	strives,
irland	irland,ireland,
hovet	court,the court,
stund	while,
östergötland	Östergötland,east gothland,
selma	selma,
amy	amy,
lady	lady,
tobak	tobacco,
strävan	the quest,
nationella	national,
skilda	separate,
miniatyr|en	thumbnail,
skilde	varied,
varandra	each other,
nationellt	national,
låga	low,
astronomer	astronomers,
inriktade	oriented,
präglades	was marked,imprinted,
stånd	position,
fönster	windows,window,
slår	switch,beats,
användbara	usable,
sålts	sold,
indikerar	indicates,
frigörelse	liberation,
berodde	depended,
agera	act,
bestämd	fixed,
strindberg	strindberg,
utskott	committee,organ,
bestämt	decided,particularly,
nsdap	nsdap,
inuti	inside,
växa	growth,grow,
kategoriledamöter	category members,category: members,
bestäms	determined,is decided,
kaffet	coffee,the coffee,
francis	francis,
drama	drama,
övertygad	confident,
ideologi	ideology,
jamaicanska	jamaican,
central	central,center,
nordliga	northernly,northern,
socialistiska	socialistic,socialist,
sri	sri,
torget	square,
bidragen	contributions,
efterkrigstiden	the post-war period,
kapten	captain,
klassiker	classic,
transporter	carriage,transports,
karriär	career,
your	your,
area	area,
sats	kit,
stark	strong,
start	start,
anställd	employed,hired,
specifika	specific,
likväl	nevertheless,still,
dopamin	dopamine,
gånger	times,
fastställa	determine,confirm,
hawking	hawking,
guillou	guillou,
wailers	wailers,
sämsta	worst,
gången	time,
traditionerna	traditions,the traditions,
expeditionen	the expidition,expedition,
minne	memory,
engelskan	english,
tidningarna	papers,
minns	remembers,remember,
miguel	miguel,
bilmärke	car make,
expeditioner	expeditions,
kostar	costs,
kungen	king,the king,
grammis	grammy,
sveriges	swedens,
godkände	approved,
styrde	steered,
knut	knut,knot,
evenemang	event,
nere	down,
drycker	beverages,
upphovsman	author,creator,
tänderna	teeh,teeth,
you	you,
köper	making,
knä	knee,knees,
drift	operation,drift,
översätts	translated,
massachusetts	massachusetts,
röda	red,
skuggan	the shadow,
tjänare	servant,
handelsmän	merchants,
morgonen	the morning,am,
färdas	travels,
susan	susan,
olympiastadion	olympa stadium,olympic stadium,
monte	assembly,
eriksson	eriksson,
beskrivningar	descriptions,
energikälla	source,energy source,energy call,
messi	messi,
öknen	the desert,desert,
loppet	bore,
antoinette	antoinette,
griffin	griffin,
råvaror	raw materials,wood,
lämpliga	suitable,
påbörjades	was started,
lämpligt	suitable,
fästning	fortress,
skiljer	differs,
vers	verse,
får	may be,can,
verk	work,works,
osv	etc.,
sanna	true,
heaven	heaven,
sverige	sweden,
behöver	need,
louis	louis,
industrialiseringen	indutrialization,industrialization,
resan	the trip,journey,
koranen	the quran,
rasism	racism,
magdalena	magdalena,
fåglarnas	the birds',birds,
egendom	property,
orgasm	orgasm,
markerade	selected,marked,
trupper	troops,
utåt	outwardly,
höja	raise,
tvskådespelare	tv actor,
besöker	visit,
bedrev	conducted,managed,
fjärde	fourth,
förbjuden	smoking,
erhöll	recieved,
bernhard	bernhard,
förbjuder	prohibiting,
misstänkta	suspected,suspect,
inblandad	mixed,
förbjudet	prohibited,
irak	iraq,
densiteten	density,
avbryta	cancel,
genomförde	carried out,
ersättare	alternate,
kronor	kronor,crowns,
observeras	observed,is noticed,
uttalat	outspoken,
lämna	leave,supply,
uttalas	pronounced,be pronounced,
arena	arena,
medarbetare	employees,
signifikant	significant,
vår	spring,
krigen	wars,
dyker	dives,shows,
stulna	stolen,
minst	at least,
boxning	boxing,
sagor	fairytales,tales,
kriget	the war,war,
hoppades	hoped,
perspektiv	perspective,
medicin	medicine,
då	then,when,
globen	lobe,
nazityskland	nazi germany,
gick	passed,
grunda	found,
dalarna	valleys,
ökat	increased,
nukleotider	nucleotides,nucleotide,
familj	family,
muslim	muslim,
avsedd	adapted,intended,
simba	pool,
arrangemang	arrangement,
taket	the roof,ceiling,
etablerad	established,
förlängningen	elongation,
planen	the plan,plan,
trummisen	the drummer,drummer,
bolagets	the corporation's,
representeras	represented,
representerar	represents,
teatrar	theaters,
massan	mass,
kurdistan	kurdistan,
reptiler	reptiles,
utökat	extended,expanded,
blodtryck	blood pressure,
latinamerikanska	latin american,
site	site,
inspelad	recorded,
räknar	counts,
räknas	calculated,are counted,
lagstiftande	legislating,
ständigt	always,constant,
mördad	murdered,murderd,
gazaremsan	the gaza strip,
ombord	onboard,board,
livslängd	life,life expectancy,
fronten	the front,
rapporterade	reported,
kejsardömet	empire,
vistelse	stay,
herrens	lord,
species	species,
gälla	valid,be valid,
serber	serbs,
ledger	ledger,
linköping	linköping,
smitta	infection,
mängden	amount,
reidars	reidars,reidar's,
ytterligare	additional,
samarbetet	co,
utför	perform,out,
long	longitude,
turkarna	turks,the turks,
torde	should,
fastän	although,
försök	experiments,
fd	former,ex,
ff	ff,
invasion	invasions,
samarbeten	cooperations,collaborations,
fn	un,the un,fn,
stabil	stable,
vattenkraft	hydroelectric power,hydro,
kostnaden	cost,
byggandet	construction,the building,
enzymer	enzymes,
allmänna	general,
korset	cross,
kognitiv	cognitive,
segrar	victories,
sänder	broadcast,transmits,
kostnader	cost,expenses,costs,
dream	dream,
nämnts	mentioned,above,
tillgångar	assets,
högst	highest,
helt	completely,totally,
bloggar	blogs,
tornet	tower,the tower,
tornen	towers,
hela	entire,full,
maffian	mafia,
hell	hell,
kombinerade	combined,
eros	eros,
hundratusentals	hundreds of thousands,
paulo	paulo,
hendrix	hendrix,
antagits	adoption,
systems	systems,
österrikes	austria's,austrias,
mahatma	mahatma,
musikalisk	musical,
bytte	swapped,
arsenal	arsenal,
konstitutionella	constitutional,
greps	was arrested,arrested,
dyrt	a high price,dearly,
petter	petter,
närmare	further,
fullt	completely,
fulla	complete,
skrivit	written,wrote,
strålning	radiation,
kontinentens	the continents,
ifk	ifk,
etnisk	ethnic,
positionen	position,the position,
märktes	labeled,
positioner	positions,
rättvisa	justice,
försäljning	sales,sale,
aktörer	players,
robert	robert,
bodde	lived,
lungorna	the lungs,
stödet	support,the support,
pythagoras	pythagoras,
känna	known,know,
efternamn	last name,lastname,
utredningen	investigation,the investigation,
heroin	heroin,heroine,
känns	felt,
delningen	pitch,
vasas	vasa,vasas,vasa's,
svarade	answered,
etnicitet	ethnicity,
skogen	woods,
skilja	seperate,separate,
american	american,
förbättrade	improved,
underhåll	support,allowance,
kung	king,
skiljs	separated,separate,
sändes	was sent,
utvecklats	developed,
synen	sight,
etiska	ehtical,
elden	fire,the fire,
riksföreståndare	regent,
minoritetsspråk	minority language,
fabriker	factories,
kallat	called,
taggar	tags,
synes	seems to,apparently,appears,
miss	miss,
rygg	back,dorsal,
deltagare	contestant,participants,
kanada	canada,
kongresspartiet	congress party,indian national congress,
station	station,
parlamentsvalet	parliament election,parliamentary elections,
nigeria	nigeria,
brittiska	british,
luminositet	luminosity,
läsa	read,
delades	divided,split,
lupus	lupus,
läst	read,
brittiskt	british,
tvungen	forced,had,
bildande	forming,formation,
växterna	plants,
brasiliens	brazil's,
långsamt	slowly,
einsteins	einsteins,
andersson	andersson,
värden	values,
värdet	the value,
stiftelsen	foundation,
gren	crotch,branch,
sekunder	second,
charlotte	charlotte,
bestämdes	was determined,
teslas	teslas,tesla's,
genomgripande	radical,good,
medeltemperaturen	the average temperature,
tvärtom	on the contrary,contrary to,vice versa,
nominerad	nominated,
militär	military,
demokratin	the democracy,democracy,
vädret	weather,
grundarna	founders,
liberalismen	the liberalism,liberalism,
lik	similar,alike,
liv	life,
mänskliga	human,
herre	lord,
avseenden	regard,
jämföras	comparable,compared,
mexiko	mexico,
åkte	relegated,
logotyp	logo,
sektor	sector,
säsongens	season,the seasons,
kan	can be,
freddie	freddie,
kap	chapter,cape,
fågel	bird,
utgör	constitutes,
himlakroppar	celestial bodies,
södra	southern,south,
förnuftet	reason,
polacker	polish,poles,
klädd	clothed,coated,
räknade	counted,
recensioner	reviews,
rådde	prevailed,was,
två	two,
osäkra	doubtful,
ingenting	nothing,
jupiters	jupiter's,jupiter,
möjligen	possibly,
counterstrike	counterstrike,
hänvisar	reference,
muslimsk	muslim,
integritet	integrity,
justice	justice,
humanistiska	humane,humanistic,
åländska	Åland swedish,aland,
ikon	icon,
lennon	lennon,
darwin	darwin,
ingå	be a part,include,be included in,
dominans	dominance,
arabvärlden	arab world,
tillhört	belonged to,
utrikes	foreign,
gått	gone,passed,
alexander	alexander,
grekiskans	greek,
restauranger	restaurants,restaurant,
avsaknaden	absence,
dömdes	sentenced,was convicted,
vilket	which,
målare	painter,
tolkiens	tolkien,
västkusten	the west coast,
grunden	base,
allmänt	generally,
maurice	maurice,
bakgrund	bakground,background,
tidigare	earlier,before,
förenta	united,
ändamål	object,purpose,
grunder	bases,
mörkare	darker,
förekom	was,
flyter	float,
direktör	director,
haddock	haddock,
pictures	pictures,
lösa	solve,
existerande	current,
pjäser	checkers,plays,
löst	solved,dissolved,1st sentence: loosely; 2nd & 3rd: solved,
läns	county,
chansen	chances,
kategorin	category,the category,
allvar	earnest,serious,
likhet	similar,resemblance,like,
utsträckning	extent,
köket	cuisine,the kitchen,
genre	genre,
länk	link,
produkter	products,
league	league,
rankning	ranking,
lejonet	the lion,lion,
anor	ancestry,
galaxer	galaxies,
boende	resident,accommodation,
viljan	will,
slavar	slaves,
kyrkliga	religious,from the church,church,
bott	lived,
läsaren	the reader,
evolutionsteorin	theory of evolution,
uppfylla	satisfy,
betydde	meant,ment,
derivata	derivative,
scientologikyrkan	the church of scientology,church of scientology,
linux	linux,
sokrates	socrates,
nacional	nacional,
skydd	protection,
merparten	most,larger part,
minskade	minimum period,was reduced,
enheten	unit,
enheter	units,
oändligt	infinity,infinitely,
konsensus	consensus,
gestalt	figure,
walter	walter,
handlingen	the story,
budgeten	budget,the budget,
anthony	anthony,
livet	the life,life,
genomfört	carried out,
genomförs	conducted,is carried out,
socialism	socialism,
hegel	hegel,
analytisk	analytical,
läser	read,are reading,
diktator	dictator,
guide	guide,
slutar	ends,end,
slutat	ended,left,
uttryckte	expressed,
nationalitet	nationality,
klippiga	rocky,
sorter	kinds,varieties,types,
bärande	wearing,leading,
lagar	laws,
tillfällen	occasion,oppertunities,
kombineras	combined,
staffan	staffan,
kombinerat	combined,
grant	word,
borgerliga	bourgeois,conservative,
deltagande	participation,
kombinerad	combined,
grand	grand,
ingår	is,
luxemburg	luxembourg,luxemburg,
folkslag	kind of people,peoples,
kungahuset	royal family,royal house,
bon	nests,
anklagats	accused,
 km	kilometers,
kommunicera	communicate,communicating,
förlag	publishers,magazine,
seglade	sailed,
armenien	armenia,
svealand	svealand,
fatta	make,to make,
kurdisk	kurdish,
stjärnorna	the stars,
präglas	characterized,
cruz	cruz,
frihetliga	libertarian,
flygplan	aircraft,airplane,
nutid	present,
präglad	marked,characterized,
innersta	innermost,inner,
feminister	feminists,
departement	department,
njurarna	the kidneys,kidney,
tortyr	torture,
skal	shell,skin,
fredliga	peaceful,
romerskkatolska	roman catholic,
uppfinnare	inventor,
kallblod	cold blooded,
filip	filip,
taiwan	taiwan,
henne	she,
gänget	the group,the gang,gang,
nikki	nikki,
barack	barack,
välkända	known,
varuhus	department store,
egenskap	trait,
djup	deep,
marco	marco,
bestå	consists,exist,comprise,
återställa	reset,
lika	similar,alike,
gör	does,makes,
kulturen	culture,
enklare	simpler,
kulturer	cultures,
gitarristen	the guitarist,
baserade	based,
unga	young,
läs	read,
immigranter	immigrants,
innan	before,
uppvärmningen	the warm-up,
känslig	susceptible,
releasedatum	release date,
dylikt	such,
infektion	infection,
gandhis	gandhi's,gandhi,
unge	kid,
donna	donna,
begärde	called,demanded,
tolkats	interpretation,interpreted,
byggnader	buildings,
biträdande	assistant,assisting,
pierre	pierre,
våldet	the violence,violence,
economic	economic,
publiceringen	the publication,publishing,publication,
syndrom	syndrome,syndrom,
sammanhängande	continous,connective,
skapat	created,
världsarvslista	world heritage list,
vilda	wild,
skapar	creates,
skapas	creates,
faktorn	factor,
slash	slash,
skapad	created,
östasien	east asia,
bägge	both,
nationalistiska	nationalistic,
sarajevo	sarajevo,
run	run,
steg	rose,
rum	room,
sten	stone,
mellankrigstiden	interwar years,
naturvetenskapliga	science,scientific,
socialister	socialists,
skrivet	written,
benfica	benfica,
bistånd	aid,assistance,
führer	fuhrer,
myndighet	authoroty,authority,
övergick	transended,went over,
linjen	line,
etablerade	established,
fysiologiska	physiological,
efterträdare	successor,
refererar	reference,
linjer	routes,lines,
edvard	edvard,
länderna	states,the countries,
ändringar	changes,
ida	ida,
egenskaper	characteristics,
ön	island,
öl	beer,
reaktorer	reactors,
institut	institution,
emellan	between,
överst	top,
föreningen	association,compound,
fokuserade	concentrated,focused,
ligga	lie,be,
spänningen	exitement,voltage,
består	exists,
visat	found,shown,
heritage	heritage,
jonsson	jonsson,
orsaker	causes,
ledamot	representative,
strukturen	the structure,structure,
japanerna	the japanese,
spektrumet	spectrum,
larry	larry,
strukturer	structures,structure,
drabbats	afflicted,
skådespelaren	actor,
skull	sake,
ute	absent,out,
nyval	re-election,election,
skuld	liability,
malin	malin,
trafikerade	frequent,trafficked,
  km²	square kilometre,
politik	politics,policies,
förbjöds	banned,forbidden,
chelsea	chelsea,
ligacupen	league cup,
bränslen	fuel,fuels,
ihåg	remember,
avsåg	meant,
sydkorea	south koreans,south korea,
hårdrock	hard rock,
igenom	through,
krigets	the war's,war,
sjunde	seventh,
musikens	music,
berättat	told,
relationerna	the relationships,
berättar	tells,
berättas	is told,
korn	korn,barley,
rester	remains,
dras	draw,preferred,
drar	earn,drag,
inkomstkälla	source of income,
william	william,
drag	characteristic,move,
mästare	master,champion,
kort	short,
resten	the rest,rest,
vindar	winds,
kors	cross,
närmaste	nearest,closest,
samarbetade	collaborated,
enade	united,
medför	entails,means,
officerare	officers,officer,
tunga	tongue,
heath	heath,
tillfälliga	temporary,
tungt	heavy,
svt	svt,
dvs	d.v.s.,i.e.,
skyskrapor	skyscrapers,
stones	stones,
bonniers	bonnier's,bonniers,
höst	autumn,fall,
placera	position,place,
indiska	indian,
katt	cat,
företeelse	feature,phenomenon,
ge	give,
tänker	thinking,
ga	ga,
go	go,
gm	by,
träd	into,tree,
kate	kate,
världsrekord	world record,
tillhör	belongs,belonging to,
toppar	tops,peak,
dröjde	not until,
sålt	sold,
wave	wave,
rinner	flow,flows,
kommunismen	communism,
försvarsminister	minister of defence,
ryan	ryan,
utbredning	distribution,distrubution,
tidszoner	time zones,
jönköping	jönköping,
stift	diocese,
akut	acute,
oklart	clear,
socialdemokratiska	socialists,social democratic,
zh	zh,
derivator	derivatives,derivative,
mussolinis	mussolini's,mussolini,
honan	the female,
geologiska	geological,
visserligen	certainly,although,
början	top,
intervjuer	interviews,
börjar	starts,starts to,start,
börjat	started,begun,
geologiskt	geologically,
svagare	weaker,
kinas	chinas,
erövringar	conquests,
hansson	hansson,
bjöd	offered,invited,
polen	poland,
bergman	bergman,
genombrott	breakthrough,
cell	cell,
experiment	experiment,
avancerade	advanced,
valen	elections,
gasen	gas,
utrikespolitiken	foreign policy,the foreign policy,
invigdes	inaugurated,
bindande	binding,
offentlig	public,published,
innerstaden	inner city,
händelsen	the occurence,event,
gåva	gift,
eminem	eminem,
vreeswijk	vreeswijk,
uppgick	was,
ryska	russian,
händelser	handelsar,events,
innebandy	floorball,
svenskans	swedish language,
västerut	west,westwards,
chans	chance,
ateism	atheism,
förening	union,compound,
kraftig	strong,
uppfinningar	inventions,
arthur	arthur,
vuxen	adult,
italienska	italian,
genetiska	genetic,
personen	person,the person,
utdöda	extinct,
genetiskt	genetically,genetic,
kunde	could,
stärka	enhance,
personer	person,people,
oktober	october,
starten	start,
nordkorea	north korea,north koreans,
invigningen	the opening,
huxley	huxley,
misslyckades	failed,
turkiets	turkey's,turkeys,
debutalbum	debut album,
microsoft	microsoft,
släppts	released,
befolkningstäthet	population density,the population density,
guds	god,god's,
kenny	kenny,
utomstående	outside,
linköpings	linköpings,
halloween	halloween,
beslöt	resolved,
studioalbum	studio album,
talat	spoken,spoke,
fördelningen	distribution,
talas	spoken,is spoken,
talar	speaks,
romantikens	romanticism,
tåget	train,the train,
kretsar	circles,circuitry,
tågen	train,the trains,
sovjetunionen	the soviet union,
fälttåg	campaign,
ferdinand	ferdinand,
folkmängd	population size,population,
kronprinsen	crown prince,the crown prince,
oroligheter	unrest,
fara	danger,
uttalet	the pronounciation,pronunciation,
dödlig	lethal,mortal,
sena	late,
fars	father,
utfördes	was carried out,preformed,
ringde	called,
österrikiska	austrian,
säljer	sells,
reagerar	react,reacts,
tillhöra	belonging to,
absint	absinthe,
encyclopedia	encyclopedia,
rörde	had something to do with,touched,was about,
kungliga	royal,
kapital	capital,
obelix	obelix,
timmar	hours,
presidenter	president,presidents,
offentliga	public,
förstördes	destroyed,was destroyed,
någonting	nothing,anything,
presidenten	president,the president,
offentligt	publicly,
verklighet	reality,
belopp	sum,
tränger	cut in,penetration,
begick	commited,
kyrkor	churches,
insekter	insects,
allting	everything,
filosofiska	philosophical,
naturgas	natural gas,
konserten	the concert,concert,
zagreb	capital of croatia,zagreb,
ägna	spend,devote,
läror	teachings,
front	front,
konserter	concerts,
dikt	poem,
intäkterna	the revenues,
miniatyr|px|den	miniature,
hunden	the dog,
kläder	clothes,
university	university,
räckte	enough,handed,
mode	fashion,mode,
förmågor	capacities,abilities,
modo	modo,
täcker	covers,
vilken	which,
föreslogs	suggested,was suggested,
illuminati	illuminati,
globe	globe,
skolgång	school attendance,schooling,
 procent	percent,per,
stiger	rises,rising,
osmanerna	ottoman turks,ottomans,
apartheid	apartheid,
skov	relapse,
skor	shoe,
sandy	sandy,
flyr	flees,
entertainment	entertainment,
förutom	except,
islamisk	islamic,
samarbetar	cooperates,collaborates,
samarbetat	collaborated,
max	max,
solsystem	solar system,
vinter	winter,
omfatta	cover,
torres	torres,
frånträde	withdrawal,
bilder	images,pictures,
lycka	happiness,good luck,
lida	sheath,suffer,
bilden	image,the image,
förstod	understood,
förbund	union,federal,
kommunala	local,municipal,
livsmedel	food,
banor	paths,line,
times	times,
åter	again,undertake,
benämnas	named,entitled,
strida	conflict,fight,
tillgången	access,
tigrar	tigers,
austin	austin,
praxis	practice,
riksdagsvalet	parliamentary election,parliamentary elections,
ursprungsbefolkningen	the native population,
minoritet	minority,
brandenburg	brandenburg,
centrum	center,
bedöma	assessment,
kategorihedersdoktorer	category of honorary degrees,
ipredlagen	ipred act,
attack	attack,
boken	paper,the book,
upphört	ceased,
dygnet	day,
infaller	no cells,falls,
final	final,
viktor	viktor,
hasch	hashish,
emellertid	however,
styrelseskick	form of government,government,
lista	list,
definierat	defined,
ben	bone,
definieras	is defined,defines,
definierar	defining,
arbetade	worked,
inbördes	relative,intermutual,
israelisk	israeli,
ber	asks,
bet	bit,
julian	julian,
kvinnans	female,
hjärna	brain,
need	need,
bordet	the table,
varade	duration,
förra	last,
tredjedelar	thirds,
visor	songs,
förlorades	lost,was lost,
släkt	family,
runorna	the runes,runes,
röst	voice,
förblev	remained,
jorge	jorge,
regn	rain,
montana	montana,
kvarstår	remains,
regi	direction,
tyskar	germans,
sändas	broadcast,be transmitted,sent,
rött	red,
planerar	planned,
skogar	forests,
långtgående	far-reaching,
platon	platon,platonic,
parker	parks,
minska	reducing,reduce,
tolkien	tolkien,
fynden	findings,
allvarliga	severe,
församling	congregation,assembly,
skedde	was,
poesi	poetry,
parken	the park,
hade	was,had,
basen	became,
baser	bases,
gemensam	common,
härskare	ruler,
förbli	remain,
varit	been,
partnern	the partner,
aspekt	aspect,
psykologin	the psyhology,psychology,
boris	boris,
klassiska	classic,
inbördeskrig	civil war,
omloppsbana	orbit,
michigan	michigan,
förbjöd	forbade,forbid,
området	the area,area,
inflytelserika	influential,
klassiskt	classical,classic,
häst	horse,equine,
områden	area,
städerna	urban,
karriären	career,the career,
älskade	loved,
gray	gray,
evolution	evolution,
processer	processes,
tillgång	access,
mohammed	mohammed,
grav	tomb,grave,
gran	spruce,
influensa	influenza,flu,
också	also,
grad	rate,
processen	the process,
vänt	turned,
produkten	product,
lätta	light,lighten,
västindien	caribbean,west india,
förband	bond,
neutralt	neutral,
landsting	county,
stats	state,
tenn	tin,
individens	the individual's,
flicka	girl,
gotiska	gothic,
staty	statue,
state	state,
företagets	the company's,
ken	ken,bank,
högra	right,
ersätta	replacing,replace,
sovjetiska	soviet,sovjet,
satsa	bet,
benämningen	the name,the designation,
merry	merry,
jobba	work,
befälet	the command,command,
problem	problems,
tjänster	services,
kaffe	coffee,
odens	odin's,node,
vulkaner	volcanos,volcanoes,
källkod	source code,
nyare	newer,
trädde	met,entered,come into effect,
varierade	varied,
älskar	loves,
stratton	stratton,
framgångsrikt	successful,
partiklar	particles,
jersey	jersey,
uppsättning	equipment,set,
fördelar	share,advantage,
helsingfors	helsingfors,helsinki,
torn	tower,
opposition	opposition,
dominerande	dominant,
kategoribrittiska	category uk,
knst	knst,
leipzig	leipzig,liepzig,
johans	johan,
revolutionen	the revolution,revolution,
johann	johann,
ovanför	above the,
kings	kings,king's,
sammanhang	connection,context,
christer	christer,
willy	willy,
trycket	pressure,
sara	sara,
fokusera	focus,
äldre	old,older,
poet	poet,
påminde	reminded,
poes	poe,poe's,
kingston	kingston,
vinci	vinci,
övertalade	persuaded,
affärer	business,
spanska	spanish,
spanien	spain,
humör	mood,
strömningar	sentiments,
kanarieöarna	canary islands,the canary islands,
 meter	meters,
erbjuda	offer,
reaktionerna	reactions,
könsorganen	the genitals,the reproductive organs,
texas	texas,
platons	plato,platos,
reaktion	reaction,
vilkas	whose,
rysslands	russia's,
enkel	simple,plain,
feber	fever,
demo	demo,removed,
rättigheter	rights,
nordirland	north ireland,northern,
måleri	painting,
kategorikrigsåret	category war years,
alfabetisk	alphabetical,
revir	turf,
reformationen	reformation,
parti	party,batch,
friidrott	athletics,track and field,
campus	campus,
varmed	whereby,
begav	traveled,
griffon	griffon,
dickens	dicken's,dickens,
korrekta	correct,
växjö	växjö,
flygbolag	airline,carriers,
anka	anka,duck,
uppnå	achieving,
nationens	nation,
rankas	ranks,
särskild	specific,particular,
införa	introducing,introduce,
eklund	eklund,
nämligen	namely,
spred	spread,
alperna	alps,the alps,
lagring	storage,
flickan	the girl,
strömmen	current,the stream,
grenar	branches,
i	in,
kärleken	love,
theodor	theodor,
lugna	calm,
europarådet	european council,
onda	evil,
rösta	vote,
störta	rush,interfere,
sänds	sends,sent,
sofia	sofia,
sofie	sofie,
förekommer	occurs,
sända	transmitting,
sände	sent,
vida	wide,broad,
jeff	jeff,
reducera	reduce,
natt	night,
nato	nato,
sweet	söt,
titta	see,
jesper	jesper,
katolska	catholic,
utan	without,
sanning	true,truth,
vanligare	more common,
historia	history,
definitivt	permanent,
historik	history,
klassificering	classification,
loss	unstuck,off,
lincoln	lincoln,
norges	norway's,
fernando	fernando,
martin	martin,
page	page,
regeringar	governments,
lager	layer,
kolonierna	colonies,
vardagliga	everyday,
pojkarna	boys,the boys,
library	library,
förlusterna	loss,
tenderar	tend,
vardagligt	everyday,
förenklat	simplified,
omöjligt	impossible,
fackföreningar	unions,
skorpan	crust,
peter	peter,
lagen	the law,
moskva	moscow,
skrifter	writings,
 km²	kilometres,
jugoslaviska	yugoslav,yugoslavian,
hyser	accomodates,holds,
folkets	the people's,people,
alliansen	the alliance,alliance,
fanns	was,
förde	out,
skriften	no.,writings,
broar	bridges,
motsättningar	oppositions,
meddelade	announced,stated,
samlades	collected,were united,
journal	journal,jurnal,
reza	reza,
kromosomer	chromosomes,
halvön	peninsula,the peninsula,
småland	småland,
usas	usa:s,u.s.,
keramik	ceramics,
freedom	freedom,frihet,
beslutade	resolved,decided,
samlats	collected,
skrev	said,
polisens	police,
troligen	likely,
hävdade	argued,claimed,
mytologi	mythology,
betydelsefulla	significant,
glenn	glenn,
underjordiska	underground,
räddade	saved,
tendenser	tendencies,
längsta	longest,maximum,
utility	utility,
hammarby	hammarby,
pc	pc,personal computer,
museum	museum,
djävulen	devil,the devil,
realiteten	de facto,reality,
afrika	africa,
distinkt	distinctive,
delstaterna	states,
instiftade	instituted,
neutral	neutral,
ho	ho,
behov	necessary,
hc	h.c.,
ha	be,
he	he,
samtida	contemporary,
svarta	black,
fysik	physics,
dator	computer,
pippin	pippin,
komiker	comic,
förslaget	the suggestion,
hästar	horses,
invandring	immigration,
bitar	bit,pieces,
farlig	dangerous,
pelle	pellet,
ordbok	dictionary,
ibland	sometimes,
erik	erik,
själ	soul,
eric	eric,
diego	diego,
omväxlande	varied,
sänktes	reduced,
moderaterna	the moderates,
speciell	specific,
mineraler	minerals,
serveras	served,is served,
vulkaniska	vulcanic,volcanic,
enastående	exceptional,
stat	state,
star	star,
liter	liters,
pontus	pontus,
revolutionära	revolutionary,
musikvideor	music videos,
stad	city,
musikvideon	music video,
resulterade	resulted,
stan	town,
bly	led,
hjärnan	the brain,
stam	tribe,
spontant	spontaneous,
etiken	ethics,
förekomma	occur,
inser	recognize,realizes,
klass	class,
alkohol	alcohol,
blogg	blog,
konsumtion	consumption,
hinner	have time to,time,
felaktig	incorrect,error,
auktoritära	authoritarian,
protest	protest,
andra	second,
fredrik	fredrik,
flest	most,the most,
buddy	buddy,
likaså	also,
upplagan	edition,
swan	swan,
kommersiellt	commercial,
kulturell	cultural,
bli	be,become,
kommersiella	commercial,
köpmän	traders,merchants,
gjordes	made,was,was made,
hemmet	the home,
kristendom	christianity,
östersjön	baltic,
vasa	vasa,
åstadkomma	provide,create,
upplysningen	the enlightenment,enlightenment,
kända	known,
kände	felt,
examen	exam,degree,
disneys	disneys,disney,
behövdes	required,
försöka	try,
chokladen	the chocolate,
avståndet	distance,the distance,
sydväst	southwest,
okänt	unknown,
sexton	sixteen,
dagens	current,todays,
upp	up,
rollfigurer	roll model,
force	force,
berlins	berlin,
förstaplatsen	first place,
bröstet	breast,
dennes	his,
avfall	waste,
neo	neo,
nej	no,
kommissionen	commission,the commission,
ned	down,bottom,
trodde	thought,
uppdelningen	division,splitting,
new	new,
representanthuset	house of representatives,
ner	bottom,
romani	romani,romany,
med	with,
genomföra	perform,out,
men	but,
drev	drove,
vinden	the wind,wind,
pedro	pedro,
mer	more,
läses	read,is read,
luther	luther,
geografiskt	geographically,
därpå	then,thereon,darpa,
tillverka	producing,
åka	go,
fyllde	filled,
ajax	ajax,
sju	seven,
kolonier	colonies,
geografiska	geographical,spatial,
dra	pulling,
snabbast	fastest,
magnusson	magnusson,
reste	travelled,
högtid	festival,
£m	million pounds,
efterföljare	following,successors,
rosenberg	rosenberg,
reagan	reagan,
inleddes	began,initiated,
fördelning	distribution,
soldat	soldier,
moral	morality,
berättelserna	the stories,stories,
datorn	pc,
gävle	gävle,
lennart	lennart,
provisoriska	provisional,
avgöra	determine,
rockband	rock band,
puls	pulse,
oscar	oscar,
ljus	light,
grundande	founding,
berlin	berlin,
anledning	reason,
wikipedias	wikipedias,
ljud	noise,
köln	köln,
kategorikvinnor	category women,
flora	flora,
trots	although,
procent	percent,
kapitalistiska	capitalistic,
sundsvall	sundsvall,
kanadas	canada's,
erövringen	conquest,
tidskriften	the magazine,magazine,
abstrakta	abstract,
världskrigets	the world war's,world war,
förväntade	expected,
talets	the speechs,
klitoris	clitoris,
konstitutionen	constitution,
tusen	thousands,
tidskrifter	periodicals,
risk	risk,
vänster	left,
satt	sat,
nobelstiftelsen	nobel foundation,
bonaparte	bonaparte,
avrättningen	execution,the execution,
trött	tired,
turnera	tour,
polis	police,
autonoma	autonomic,
stilla	still,stationary,
tycktes	seemed,
orsakar	causes,
orsakas	caused,causes,
orsakat	caused,
utomeuropeiska	overseas,non-european,
gård	farm,house,
könsorgan	sex organ,
klarar	do,
president	president,
orsakad	caused,induced,
indelat	divided,split,
medföra	result,
indelas	divided,
indelad	divided,
medfört	resulted,led to,
låtskrivare	songwriter,
självklart	course,
indisk	indian,
ändra	change,
kvicksilver	mercury,witty zeal,
förfäder	ancestors,
fifa	fifa,
föreställningen	the concept,show,
panthera	panthera,
ibrahimović	ibrahimovic,
munnen	the mouth,mouth,
murray	murray,
föreställningar	performances,
helena	helena,
buddhister	budhists,buddhists,
listor	lists,
personal	personal,staff,
förödande	devastating,
amerikanen	american,
amerikaner	american,
irans	iran's,
federationen	federation,
friska	fresh,
aborter	abortions,
infektioner	infections,infection,
startar	begins,start,
downs	down,
stimulerar	stimulating,
miljon	million,
myntades	coined,was coined,
huvudrollen	leading part,the main role,
inledde	started,launched,
tillvaron	life,
sida	page,side,
överraskande	surprisingly,
skeppet	nave,
side	side,
kammaren	chamber,the chamber,
liga	compatible,league,
päls	fur,
mediet	medium,
medier	media,
milan	milan,
aids	aids,
håret	hair,the hair,
kiev	kiev,
uppsala	uppsala,
årsåldern	years old,
hänvisa	reference,refer,
talet	rate,
ihop	up,together,
talen	rate,years,
sluta	end,stop,
återfanns	was rediscovered,found,
venezuela	venezuela,
bestod	was,
foto	photo,
neutroner	neutrons,neutron,
larssons	larsson's,
normer	standards,
stöds	is supported,
nietzsche	nietzsche,
nomineringar	nominations,
uppförande	code,behavior,
folkvalda	elected,
faktum	fact,
iso	iso,
reinfeldt	reinfeld,
representant	representative,
sökte	searched,
starta	start,launch,
stewart	stewart,
gå	go,
nätet	net,
jordanien	jordan,
arrangeras	arranged,
skalvet	quake,
leddes	was led,
massiv	massive,
objektet	object,
föreslagit	suggested,
girls	girls,
vikingatiden	the viking age,vikings,
förbi	past,
objekten	the objects,
hollywood	hollywood,
någonstans	somewhere,nowhere,
alfred	alfred,
åskådare	spectators,
medeltiden	middle ages,
besegrades	defeated,
skaffade	acquired,aquired,
sabbath	sabbath,
grönwall	gronwall,
symptom	symptoms,
hundar	dogs,
chef	head,
formell	formal,
kontrast	contrast,
antarktis	antarctica,antarctic,
street	street,
regissören	director,
härkomst	origin,
parter	sides,
troligtvis	probably,
bobo	bobo,
palace	palace,
stadsdelen	the district,district,
låta	let,
mina	my,mine,
modern	modern,
självständiga	independent,
självständigt	independent,independently,
triangel	triangle,
tecken	sign,
lämnar	leaves,
lämnas	left,
lämnat	left,
skildringar	descriptions,
tidiga	early,
monetära	monetary,
muskler	muscles,
italiens	italy's,
tidigt	early,
tål	is resistant to,
blue	blue,
dessa	these,
bildar	serves as,form,
bildas	formed,
tåg	rail,trains,
bildat	formed,
dödsfall	deaths,
luthers	luthers,
verksamma	active,
marie	marie,
typ	type,
diskuterats	been discussed,discussed,
maria	maria,
don	don,
dom	conviction,
materiella	material,
härstammar	derived,stems,
slipknot	slipknot,
läsare	readers,reader,
points	point,
följande	following,the following,
dos	dosage,
kristen	christian,
långvariga	long,long-standing,
koppla	coupling,
införde	introduced,
hjälper	helps,shows,
västeuropa	western europe,
befälhavare	commander,
liza	liza,
droger	drugs,
skyldig	responsible,guilty,
långvarigt	prolonged,long-standing,
nevada	nevada,
odling	cultivation,
krönika	chronicle,
anländer	arrives,
helhet	whole,
monica	monica,
stycke	piece,
meningar	sentences,
kollapsade	collapsed,
stop	stop,
stor	large,
stol	chair,seat,
präster	priests,
christopher	christopher,
stod	stood,
mönster	marks,
earl	earl,
bar	bar,
bas	base,
skrivas	printed,
existerat	existed,
anlades	was built,
fokus	focus,
förändra	change,
gärningar	deeds,
anknytning	tie,
zonen	the zone,
zoner	zones,
gunnar	gunnar,
dittills	thus far,so far,
vände	reversed,
turnén	turn,
öppnade	opened,opening,
inledningsvis	by way of introduction,
skrevs	was,
naturligtvis	course,naturally,
skrift	no.,
underart	subspecies,
sorts	variety,
göta	göta,
omkringliggande	surrounding,
smguld	sm gold,gold medal in the swedish championships,
artikel	article,
armeniska	armenian,
kämpa	fight,
motto	motto,
typisk	typical,
isotoper	isotopes,
fns	un's,tris,
regering	the government,government,
näringslivet	business,industrial life,
fördraget	the treaty,treaty,
fördragen	treaties,the compacts,
kol	charcoal,
ung	young,
ernst	ernst,
regelbunden	regular,
obamas	obama,obama's,
atombomberna	the nuclear bombs,
mellanrum	space,gap,
nationalförsamlingen	national assembly,
synsättet	view,
avsikt	intends,
interna	internal,
omstritt	controversial,
varmt	hot,
basis	basis,
sidan	side,
kallats	called,
blodkroppar	blood cells,
cyrus	cyrus,
varma	hot,
frisk	healthy,fresh,
tillämpa	administer,applying,
idol	idol,
betydelsefull	meningful,
igång	start,start up,
provinsen	province,
utseende	appearance,
sällskapshundar	pet dogs,companion dog,
namnen	names,name,
mindre	smaller,less,
etniskt	ethnic,
azerbajdzjan	azerbaijani,
etniska	ethnic,
pornografi	pornography,
ix	the ninth,
förgäves	in vain,
albaner	albanians,
mexico	mexico,
kvinnor	female,
ip	ip,
sushi	sushi,
it	it,
hämnd	revenge,
ik	ik,
huvudort	main town,principal town,
im	im,
il	il,
in	in,
colosseum	colosseum,
utgåva	edition,
stoppa	stop,
konkurrensen	the competition,competitive,
vänstern	western,
make	make,husband,
producerats	produced,
bella	bella,
västberlin	west berlin,
kommunistpartiets	communist party,the communist partys,the communist party,
roland	roland,
därmed	therefore,
industriell	industrial,
makt	power,
benämningar	terms,
anglosaxiska	anglo-saxon,
atmosfären	atmosphere,the atmosphere,
skickades	was sent,sent,
kim	kim,
nicklas	nicklas,
folkrikaste	populous,most populus,
akademiska	academic,
protesterna	the protests,
roms	romes,roms,
vetenskaplig	scientific,
sydamerika	south america,
dåvarande	then,formerly,
värmland	wermlandia,värmland,
roma	roma,
viktiga	important,
grannländer	neighbors,neighboring countries,
facto	facto,
just	right,just,
kongressen	congress,
jämför	compare,
sporting	sporting,
universitet	university,
psykos	phychosis,psychosis,
bollen	the ball,
västeuropeiska	western european,
zon	zone,
human	human,
anders	anders,
beskriver	describes,
premiärminister	prime minister,
fysiker	physicist,
hävdar	states,assert,
bokstäver	letters,
troligt	likely,
hävdat	argued,claimed,
självstyrande	self-governing,independent,self-governance,
strax	soon,just,
royal	royal,
julen	julien,christmas,
jules	jules,
friedrich	friedrich,
amerikas	america,
massa	mass,
borgen	castle,bail,the castle,
komintern	comintern,
språkets	the language's,language,
arkitekturen	the architecture,
gustav	gustav,
behövde	did,
särdrag	features,
följaktligen	consequently,
författningen	constitution,
bekräftar	confirmed,
gustaf	gustaf,
trafikeras	served,trafficked,
trafikerar	traffic,frequent,
bekräftat	confirmed,
världsdel	continent,
medborgarskap	citizenship,
kommunerna	kommunera,the municipalities,
släkting	relative,
intensiv	intensity,
litauen	lithuania,
syrien	syria,
kemiska	chemical,
vattnet	the water,
kontinent	continent,
kunna	to,be able,
dead	dead,
befolkningen	the population,population,
uppmärksammades	attention,drew attention,
jupiter	jupiter,
befann	located,
kemiskt	chemically,
statistik	statistics,
oralsex	oral sex,
kommuner	municipalities,local,
hudfärg	color,
miljöproblem	environmental problem,environmental problems,
normal	normal,
hittar	found,finds,
däggdjuren	mammals,the mammals,
säsongerna	seasons,
shakespeare	shakespeare,
hertig	duke,
filmatiserats	cinematized,been filmed,
benämns	designated,is mentioned,
knep	tricks,
angrepp	attack,
burj	burj,
versioner	versions,
bolt	bolt,
härstamma	stem,
burr	burr,
förkortas	reduced,
förkortat	shortened,abbreviated,
irländska	irish,
flyttat	moved,
fördelen	advantage,the advantage,
ljungström	ljungstrom,ljungström,
därutöver	addition,moreover,
maskiner	equipment,
omröstning	vote,
mycket	very,much,
tillverkas	manufacture,
magazine	magazine,
ishockey	ice hockey,hockey,
strömmar	streams,flow,
grenen	the branch,branch,
förknippade	associated,
äktenskap	marriage,
psykisk	psychic,mental,
français	francais,
grundades	founded,was founded,
jens	jens,
romulus	romulus,
orsak	factor,
spåra	track,
amsterdam	amsterdam,
havsnivån	sea level,
fastlandet	mainland,
estniska	estonian,
märks	labeled,noted,
tennis	tennis,
könen	the sexes,
bönder	farmers,
bolivia	bolivia,
märke	label,
hyllade	acclaimed,
själv	alone,own,himself,
ford	ford,
berg	mountain,
japansk	japanese,
bero	depend,due,
bättre	better,
epoken	epoch,the epoch,
fort	fast,quickly,
definierade	defined,
spelade	played,
positiv	positive,
slaviska	slavic,
flickvän	girlfriend,
regeringen	the government,
båten	vessel,the boat,boat,
skelett	skeleton,
månens	the moon's,the moons,
avsnitt	section,part,episode,
phil	phil,
försörjde	living,
uttryckligen	specifically,
handelspartner	trading partner,
tosh	tosh,
kanske	may,
primtal	prime number,
byggnaden	building,the building,
vista	vista,
handen	hand,
handel	trade,
kunnat	could have been,
svärd	sword,
digital	digital,
betalt	charge,
marxism	marxism,
kungamakten	monarchy,the monarchy,
sades	was said,
överenskommelse	deal,arrangement,
frodo	frodo,
exporten	the export,
katekes	catechism,
accepterade	accepted,
engagemang	commitment,
riktad	directed,
ökande	increasing,rising,
fss	fss,
expandera	expand,
riktat	directed,pointed,
riktas	direct,target,
riktar	targets,target,
armar	arms,
bomben	the bomb,
telefon	telephone,
spår	track,
manager	manager,
bomber	bombs,
vikingarna	the vikings,
marissa	marissa,
dä	the elder,
imperiet	the empire,empire,
avbrott	break,breaks,
uppdelning	partitioning,
petersburg	petersburg,
dö	die,
me	me,
illa	bad,
din	your,
die	die,
dig	up,
trenden	the trend,
afrikansk	african,
höjdes	increased,was raised,
dit	there,where,
spets	tip,point,
bulgarien	bulgaria,
olympia	olympia,
ville	did,wanted,
malmö	malmö,malmo,
diskografi	discography,
villa	house,villa,
slagit	held,
reklamen	the commercial,advertising,
invandringen	immigration,
rymden	space,
utlösning	release,ejaculation,trigger,
hästen	the horse,
bakom	behind,
afghanistan	afghanistan,
viktig	major,important,
kokain	cocaine,
föredrog	preferred,
lönneberga	lönneberga,lonneberga,
somalia	somalia,
international	international,
madagaskar	madagascar,
nationalismen	nationalism,
tibet	tibet,
henry	henry,
högkvarter	headquarters,head quarter,
avsaknad	absence,
kommun	local,municipality,
beskrivits	described,
boy	boy,
diagnoser	diagnoses,
canadian	canadian,
bor	lives,
gyllene	golden,
folkmun	colloquially,
bok	book,
mängder	amount,
extrem	extreme,
mänsklighetens	humanity's,humanities,
bolivianska	bolivian,
diagnosen	diagnosis,the diagnose,
hotell	hotel,
sporter	sports,
enorma	enormous,
utövar	carrying,exercise,
utövas	is practised,exerted,exercised,
världshälsoorganisationen	world health organization,
asiatiska	asian,
sporten	the sport,port,
religionsfrihet	religion,religious freedom,
enormt	gigantic,fusionenormously,
platån	sycamore,the plateau,
skräck	horror,fear,
hemmaarena	home ground,
tennisspelare	tennis player,
semifinalen	semi finals,
peru	peru,
kristian	kristian,
statsmakten	the government,power,
österrikeungern	oster kingdom hungary,austria-hungary,
detaljer	details,
avsattes	dismissed,
brukade	used to,
ögon	eyes,
kemisk	chemical,
fly	escape,
hända	may,
hände	happened,
tokyo	tokyo,
mästarna	the champions,
söka	search,searching,
träffades	met,was met,
vittnen	witnesses,
akademien	the academy,academy,
präglade	characterized,
anslutna	connected,
bristande	wanting,lack,
sökt	pending,
ulf	ulf,
hiroshima	hiroshima,
kenneth	kenneth,
uruguay	uruguay,
winston	winston,
agent	agent,
bemärkelse	meaning,sense,
skadades	was wounded,damaged,
council	council,
dennis	dennis,
kunglig	royal,
diskuterades	discussed,
oslo	oslo,
engelsmännen	the english,the british,
återvänder	returns,
varor	products,
ekonomiska	economic,economical,
till	to,
gitarrist	guitarist,
nya	new,
nye	new,
regeringstid	term of government,
överensstämmer	conform,agree,
uppföljare	sequel,
fotboll	football,
läkare	doctors,doctor,
maj	may,
mao	mao,
man	is,one,
asien	asia,
johnson	johnson,
kulturella	cultural,
sådana	such,
eng	eng.,
tala	speaking,speak,
block	block,
basket	basketball,
romantiken	romance,romanticism,
nå	access,
sådant	such,
lsd	lsd,
bussar	bus,
bevisa	prove,
alfabetet	alphabet,the alphabet,
unionen	the union,
gällde	applied,applied to,was,
sällsynta	rare,
moralisk	moral,
huvudsak	main thing,
lyrik	poetry,
motståndet	the resistance,the resistence,
verksam	active,
landskap	province,landscape,
juryn	jury,
sekter	sects,
äkta	married,genuine,
nazisterna	nazis,
policy	policy,
växte	grew,
main	main,
utgjorde	made up,was,
lägst	lowest,
steget	step,
kräver	requires,
janeiro	janeiro,
domstolar	courts,
försörjning	sustentation,supply,
sibirien	siberia,
leds	passed,
vindkraft	wind power,
färg	colors,colour,
uppskattning	appreciation,estimated,
leda	lead,
villkoren	the terms,conditions,
rock	rock,
föremål	object,subject,
tysklands	germany's,germanys,
guevara	guevara,
latin	latin,
tacitus	tacitus,
hellre	more preferably,rather,
söner	sons,
vattendrag	streams,watercourse,
avkomma	progeny,offspring,
girl	girl,
saudiarabien	saudi arabia,
canada	canada,
jackson	jackson,
håkansson	hakansson,håkansson,
avrättningar	execution,
pamela	pamela,
områdena	the areas,
tronföljare	heir apparent,successor,
kattdjur	felidae,cat,
premiären	premiere,
ansiktet	face,
monster	monsters,
ort	neighborhood,location,
konstnär	artist,
chiles	chiles,chile's,
oro	anxiety,
dubbla	double,
california	california,
miley	miley,
kognitiva	cognitive,
ord	word,
tunnelbanan	the subway,metro,
gott	good,
upplevde	experienced,felt,
preventivmedel	contraceptives,
självmord	self-killing,suicide,
uppvisar	shows,
rankningar	rankings,
vision	vision,
stängdes	closed,
first	first,
centrala	central,
grupperna	groups,
intryck	appearance,
uttalanden	statements,
här	here,
rachel	rachel,
folklig	folk,
lat	methacrylate,
centralt	central,centrally,
skapandet	creation,the making,
kommunism	communism,
grundämnet	the element,
missnöje	dissatisfaction,
homogen	homogenous,
visar	is,shows,
visas	shown,
västbanken	the west bank,
grundämnen	elements,
individ	individual,
örebro	Örebro,
öronen	lugs,the ears,
besluten	decisions,
anus	ass,anus,
köpenhamns	copenhagen,copenhagen's,
fysiska	natural,physical,
fysiskt	physical,
danny	danny,
löstes	solved,dissolved,
drevs	concentrated,was driven,
beslutet	the decision,
konkreta	specific,
fiender	enemies,
fienden	enemy,the enemy,
medlemmarna	the members,
lugn	calm,
jordytan	earth crust,
fordon	vehicle,
inträde	entry,
marklund	marklund,
jämlikhet	equality,
stadsdelar	districts,city districts,neighborhoods,
marijuana	marijuana,
större	greater,bigger,
formerna	forms,
tänder	teeth,
orsakerna	the causes,
kevin	kevin,
adeln	nobility,
nikola	nikola,
politiska	political,
förälskad	in love,
menas	mean,
skulptur	sculpture,
centralbanken	central bank,
politiskt	political,
performance	performance,uppträdande,
centralstation	central station,
channel	channel,
riktningar	direction,
norman	norman,
teoretiska	theoretical,
morden	murders,
dagbladet	dagbladet,
halvan	half,
politisk	political,
teoretiskt	theoretic,theoretical,
mordet	murder,
arbetat	worked,
civilisationer	civilizations,
otaliga	countless,
lojalitet	loyalty,
drottning	queen,
grammatik	grammar,
österut	eastwards,
kontrolleras	is controlled,controlled,
kontrollerar	controls,
ungdom	youth,
civilisationen	civilization,
show	show,
adolfs	adolf's,adolf,
regioner	regions,
generalsekreterare	the secretary-general,secretary general,
samlingsalbum	compilations,
helig	holy,
dick	dick,
historier	stories,
passande	fitting,suitable,matching,
historien	history,
black	black,
medeltidens	medieval,
experimenterade	experimented,
ges	be given,
ger	give,gives,
raser	races,
klasser	classes,
kulturellt	culture,cultural,
konsolen	bracket,
motsvarande	corresponding,
skådespelare	actor,
inspelningarna	recordings,
personliga	personal,
vintergatan	milky way,the milky way,
firade	celebrated,
ledaren	conductor,
gen	gene,
beskyddare	protector,patron,
himmlers	himmlers,
mattis	mattis,
bengtsson	bengtsson,
statistiska	statistical,
dianno	di'anno,dianno,
spridda	spread,
europacupen	european cup,
london	london,
tolfte	twelth,twelfth,
relativt	relative,relatively,
sämre	poor,
sekulära	secular,
fokuserar	focuses,focus,
toppade	topped,
relativa	relative,
sean	seab,sean,
slöt	closed,
utgiven	published,
menat	meant,
menar	means,
kandidater	candidates,
försvarsmakten	national defense,
visades	was,
vanns	was won,
personligt	personal,private,
erövrades	conquered,concoured,
människas	human,
landets	the country's,its,
tsaren	the czar,czar,
august	august,
ju	the,
forskaren	researcher,
jr	jr.,junior,
åker	go,
timme	hour,
tum	inch,
fick	was,
signaler	signals,
lexikon	lexicon,
kirsten	kirsten,kristen,
ministrar	ministers,
rugby	american fotboll,rugby,
ån	from,the river,
utvalda	selected,
tour	tour,
paret	pair,the couple,
ås	ridge,
år	the year,year,
vätska	liquid,
tryck	press,print,
väst	west,the west,
århundraden	centuries,
cancer	cancer,
statschefen	the head of state,
syntes	synthesis,
grundare	founder,
territorium	state,
mätningar	measurements,measurments,
ryggen	the back,back,
barry	barry,
överföra	transmit,transfer,
bildats	formed,
ja	yes,
västliga	western,
utsatta	exposed,
mars	march,
överförs	is transferred,
plötsligt	suddenly,
marx	marx,
mary	mary,
kultur	culture,
nederländerna	the netherlands,netherlands,
flaggan	flag,
cobain	cobain,
partido	partido,
avskaffa	abolish,
bmi	bmi,
jagar	hunting,
spelfilmer	motion pictures,feature film,feature films,
klädsel	cover,
meningen	sense,
fortsatt	further,continued,
metall	metal,
dragit	dragged,preferred,
uppstod	developed,was,
kategorimän	category: men,category men,
insåg	realized,
nionde	ninth,
sahara	sahara,
intressanta	interesting,
uppmanade	urged,
liknande	similiar,similar,
uppfyller	fulfills,
hålls	maintained,is held,
par	pair,
jesu	jesu,
edwin	edwin,
lava	lava,
hålla	hold,keep,
röka	smoking,
stött	met,supported,
pan	pan,
samt	also,as well as,
tidvis	times,
hösten	fall,the fall,the autumn,
kuba	cuba,
teknisk	technical,
lösningar	solutions,
sömn	sleep,
fattas	taken,
bang	bang,
wahlgren	wahlgren,
identifiera	identification,
gates	gates,
münchen	munich,
bebyggelse	settlement,settlements,
privatliv	private,
reaktionen	reaction,
dinosaurierna	dinasaurs,
skapelse	creation,
vilja	will,like,
byggnad	building,
reaktioner	reactions,
våld	violence,force,
jakten	the hunt,hunt,
ideologiskt	ideological,
grannländerna	neighbors,
bowie	bowie,
avskaffandet	abolishment,
gotland	gotland,
ideologiska	ideological,
motverka	counteract,
trä	wood,
möter	meets,
vintern	the winter,winter,
schwarzenegger	schwarzenegger,
underarten	subspecies,
mån	concerned,
mor	mother,
haft	had,
prägel	character,mark,
tillbehör	accessory,
kategori	category,
jakt	hunt,hunting,
temperatur	temperature,
mon	mon,
underarter	subspecies,
baltiska	baltic,
kollektiv	collective,public,
mod	courage,
christina	christina,
adams	adams,
födda	born,
började	started,began,
födde	gave birth too,born,
jordbävningar	earthquakes,
manhattan	manhattan,
mänsklig	human,
sågs	observed,was observed,
göran	göran,
bipolära	bipolar,
göras	be made,
rikskansler	chancellor,
kategorisveriges	category sweden,
feodala	feudal,
maos	maos,mao's,
förs	led,out,
jordbruket	the agriculture,
lotta	raffle,
fört	lead,
reportrar	reporters,
föra	pre,
ända	as far as,up,
demokratisk	democratic,
traditionell	traditional,conventional,
samman	together,
moderata	moderate,
vistas	present,
tunnlar	tunnels,
londons	london's,
cellen	cell,the cell,
olof	olof,
akon	akon,
sjätte	sixth,
celler	cells,
förhistoria	prehistory,
island	icelandic,
allians	alliance,
metaforer	metaphores,
lands	land,on land,
lagarna	the laws,
retoriken	rhetoric,
herbert	herbert,
matematiska	mathematical,
arvid	arvid,
wilde	wilde,
beskrivas	described,be described,
einstein	einstein,
mark	ground,
intellektuella	intellectuals,intellectual,
floderna	floods,rivers,
fullständigt	full,
gravid	pregnant,
behandling	treatment,
varelse	creature,
emellanåt	once in a while,occasionally,
anfalla	attack,
välmående	healthy,prosperous,
fullständiga	full,complete,
kvinnlig	females,female,
tillfälligt	temporarly,temporary,
eget	own,
utbredd	widespread,spread,
härifrån	from here,here,
e	e,
egen	own,
tävlingen	competition,contest,
vhs	vhs,
exemplar	copies,example,
bibliografi	bibliography,
manuel	manual,
verkliga	fair,
identifierade	identified,
humanismen	humanism,
parlament	parliament,
håkan	håkan,
följde	followed,
youtube	youtube,
öns	the islands,
prestigefyllda	prestigious,
skriven	written,
palats	palace,
arabiska	arabic,arabian,
goebbels	goebbels,geobbels,
film	film,
again	again,
genrer	genres,
vanliga	regular,usual,
istanbul	istanbul,
spåren	the tracks,wake,
rubiks	rubiks,rubik's,
muren	wall,
produktiv	productive,productivity,
stannade	stayed,
spåret	groove,
genren	genre,
faktorer	factors,
däremot	on the contrary,
ordna	arranging,arrange,
profet	prophet,
ungarna	kids,the young,
förändrade	changed,
rykten	rumors,
ledning	conduit,guidance,
henriks	henry,
kyros	cyrus,
chris	chris,
medicinska	medical,
dvärghundar	miniature dogs,
nöjd	content,
palestinska	palestinian,
uppfostran	upbringing,
medicinskt	medical,
god	good,
snabbaste	fastest,
begå	commit,
resolution	resolution,
åtskilda	separated,separate,
mellanöstern	middle,the middle east,
vila	rest,
socialismen	socialism,
dollar	dollar,
vill	to,
hindrar	prevent,prevents,
ingripande	negative,
inspirerad	inspired,
liam	liam,
levern	the liver,liver,
zink	zinc,
symbolen	the symbol,
kategorilevande	category of live,
rwanda	rwanda,
symboler	symbols,
skydda	protection,
skriver	type,
seriens	series,
kasta	discard,throw,
avhandling	thesis,
israeliska	isrealic,
fall	where,
ramen	frame,
behöva	need,
kulminerade	culminated,
miljoner	millions,
båtar	boats,
bröderna	brothers,the brothers,
suttit	been,sat,
ockuperades	occupied,
cornelis	cornelis,
massor	lots,tons,
växthuseffekten	the greenhouse effect,
intressant	of interest,
material	material,materials,
abc	abc,
danmark	denmark,
abu	abu,
public	public,
lärare	teacher,
långhårig	long haired,
bebott	inhabited,
närhet	close,closeness,
legat	formed,
jonas	jonas,
free	free,
benen	legs,
valt	chosen,selected,
sångare	singer,
historiker	historians,
jackie	jackie,
faktiskt	actually,
uppslagsverk	encyclopedia,
alexandria	alexandria,
sjukhuset	hospital,
africa	africa,
nacka	nacka,
släktingar	relatives,
varianterna	variants,the diversities,
rösterna	votes,
författaren	the author,author,
hyllning	tribute,
eye	eye,
medlem	member,
torrt	dry,
utmärkelsen	award,the award,
utmärkelser	awards,
torra	dry,
diamond	diamond,
människa	human,man,
romersk	roman,
koma	coma,
tillkommer	reside,will be,
hundraser	breed of dogs,breeds,
skivor	plates,records,
vladimir	vladimir,
länkar	links,
des	des,
det	is,
roosevelt	roosevelt,
del	part,
lindgren	lindgren,
den	it,
befintliga	current,existing,
samtliga	all,
hastigt	rapidly,fast,
latinets	latin,the latin,
sovjetunionens	soviet union,
betoning	stress,
hjälpte	helped,
sjukdom	illness,
medförde	resulted,brought,
födseln	birth,the birth,
sträng	string,
robinson	robinson,
protein	protein,
makten	power,the power,
hämta	retrieve,fetch,
stil	type,
psykotiska	psychotic,
georgien	georgia,
stig	stig,
verkligheten	real,reality,
blad	leaves,
försvinner	disappears,
primära	primary,
vikten	importance,weight,
makter	powers,
hoppade	jumped,
avtalet	the contract,
pettersson	pettersson,
laboratorium	laboratory,
ännu	even,yet,
judiska	jewish,
huvudkontor	central office,headquarters,
ligger	is,
vatten	water,
rastafarianer	rastafarian,
rockgrupper	rock bands,
facebook	facebook,
paz	paz,
konservatismen	conservatism,
civila	civil,
inåt	inwards,inwardly,
nordsjön	north sea,
officiella	official,
latinamerika	latin america,
fältet	the field,field,
höll	gave,
göra	do,
mörkt	dark,
gradvis	gradually,progressively,
tvåa	second,
baltikum	the baltics,baltics,
mörka	dark,
görs	is,is made to,
officiellt	official,officially,
människans	humans,mankinds,human,
längden	lenght,
diskussion	discussion,
ärftliga	genetic,
edmund	edmund,
inbördeskriget	civil war,
andré	andre,
odlade	grew,cultured,
saknades	missing,
trossamfund	religious communities,
suverän	terrific,sovereign,
good	good,
träffar	meets,hits,
ställas	set,be set,prepared,
planerna	the plans,
fängelse	prison,
sexuellt	sexual,
oxford	oxford,
skrifterna	scriptures,
association	association,
toronto	toronto,
robbie	bobbie,robbie,
kungarna	the kings,kings,
namibia	namibia,
out	out,
byggt	building,built,
anslöt	joined,
trådlös	wireless,
fisk	fish,
energy	energy,
hard	hard,
flytta	move,
byggs	building,
förenade	united,
energi	energy,
seder	subsequently,custom,
perry	perry,
sanningen	truth,the truth,
östman	Östman,
sällsynt	rare,
oftast	usually,most often,
infrastrukturen	infrastructure,
ölet	the beer,beer,
forskning	research,
perro	perro,
förföljelser	pursuits,persecutions,
fullständig	full,complete,
konflikt	conflict,
prins	prince,
lawrence	lawrence,
strömning	flow,
blekinge	blekinge,
uralbergen	urals,
eventuellt	eventually,
viken	gulf,
helsingör	elsinore,helsingör,
inflationen	inflation,
investeringar	investments,
finland	finland,
jordens	earth,
utöver	addition,
fått	was given,with,
styre	governance,rule,
legenden	legend,
ensam	alone,
styra	controlling,steer,
top	top,
sjunkande	decreasing,
dont	do,
säkerhetsråd	security,security council,
treenighetsläran	doctrine of the holy trinity,trinity,school of trinity,
snarast	rather,as soon as possible,
juridiska	legal,
carter	carter,
förklarade	explained,said,
kom	came,
diskriminering	discrimination,
kon	group,
noga	carefully,
observationer	observations,
förhindrar	prevents,prevent,
kategoriasiens	category of asia,
kardinal	cardinal,
järnvägar	failways,rail,
triangeln	triangle,the triangle,
part	party,
gudarna	the gods,
domstolen	court,the court,
direkta	direct,
matteusevangeliet	gospel of matthew,
följden	result,
b	b,
avtal	agreement,contract,
proteinerna	proteins,
dogs	dogs,
personens	person,the persons,
singapores	singapores,
hellström	hellström,
baháí	baha'i,bahá'í,
avtar	declines,avatar,
självständig	independently,
följder	impact,
följdes	followed,was followed,
rikedom	riches,
försökte	try,tried,
bränsle	fuel,
gjord	made,
flertalet	most,
gjort	made,done,
mountain	mountain,
hundratals	hundreds of,hundreds,
mussolini	mossolini,
infrastruktur	infrastructure,
caesar	caesar,
genast	at once,immediately,
taktik	strategy,
dramatiskt	dramatically,
skjuta	delay,
militärt	military,
patterson	patterson,
krafter	forces,
gillade	liked,
niclas	niclas,
kraften	the force,
utbrott	outbreak,
samtidigt	while,
organiserade	organized,
högt	high,highly,
ko	co,cow,
km	km,kilometers,
kl	at,
kr	kronas,
liechtenstein	liechtenstein,
organisk	organic,
thomas	thomas,
venedig	venice,venedig,
kvalitet	quality,
byttes	was exchanged,
relation	ratio,relation,
utveckla	developing,
fina	beautiful,fine,
nämns	mentioned,
antagit	adopted,presumed,
konto	account,sign,
undre	lower,
wallenberg	wallenberg,
medverka	take part,participate,
världens	the world,the worlds,
tionde	tenth,
religionerna	religions,
förbudet	ban,the union,
avseende	regard,for,
blomstrade	flourished,
typiskt	typically,typical,
nationalpark	national park,
notation	notation,
beslutar	decides,
vänskap	friendship,
express	express,
beslutat	resolved,
förklarat	explained,declare,
typiska	typical,
förklarar	explains,
gamla	ancient,old,
husen	housing,the houses,
skickas	is sent,
skickar	sends,
brukar	usually,
wallander	wallander,
gamle	old,
uttrycket	the expression,expression,
uttrycker	expressing,
flykt	escape,
huset	housing,
svarar	responds,
somrar	summers,
stadium	stage,
styrdes	governed,
suveränitet	sovereignty,
rollfigur	character,
godkännas	approved,be approved,
höglandet	the highland,
tengil	tengil,
rovdjur	predator,
fans	fans,
landsbygden	rural,rural area,
champagne	champagne,
romarriket	roman empire,the roman empire,
bildandet	formation,establishment,
professionella	professional,
framförs	is presented,performed,
framfört	expressed,
rörelserna	the movements,movement,
kritiserades	critisized,
framföra	express,convey,
marilyn	marilyn,
musklerna	muscles,the muscles,
statligt	state,governmental,
uppfattning	understanding,view,
praktiskt	convenient,
statliga	state,
restaurang	restaurang,restaurant,
romska	romani,roma,
beta	graze,beta,
globala	global,
kroatiens	croatias,
förklaring	explanation,statement,
folkmord	genocide,
karaktären	character,
andas	breathes,
karaktärer	characters,
således	hence,thus,
tennessee	tennessee,
globalt	globally,global,
behöll	kept,retained,
försäljningen	sales,
lyfta	lift,
våningar	floors,storeys,
laos	laos,
bestämde	chose,
inför	before,
bengt	bengt,
popularitet	popularity,
gav	gave,
effektiva	effective,
gas	gas,
vana	familiar,
kalmar	kalmar,
effektivt	effective,
trupperna	troops,the troops,
detsamma	the same,
bild	image,
motorväg	freeway,highway,
åtalades	was charged,was prosecuted,
spridning	diffusion,distribution,proliferation,
bill	car,
döptes	baptised,
portugal	portugal,
arenan	arena,
påbörjade	started,
monroe	monroe - it's a persons name,monroe,
rederiet	the shipping company,shipping company,
dödat	killed,
granska	examining,
sjuk	disease,
dödar	kill,kills,
dödas	killed,
hamna	end,
motståndaren	the opponent,opponent,
administrationen	administration,
dödad	killed,
tyder	indicates,
sapiens	sapiens,
övertogs	were taken,overtaken,
skotska	scottish,
syd	south,
jerusalems	jerusalem's,
moment	step,
kallades	was called,called,summoned,
parentes	brackets,
avsett	avset,intended,
nämnde	mentioned,said,
mot	against,
nämnda	said,
kungariket	kingdom,
noll	zero,
kapitel	chapter,
albanien	albania,
jorderosion	earth erosion,soil erosion,
ministerrådet	minister counsellor,
skott	shots,
albanska	albanian,
norrland	norrland,northern,
dikter	poems,
bibeln	bible,
kommunister	communists,
juventus	juventus,
organization	organization,
representanter	representatives,
passerar	passes,pass,
struktur	structure,
senaste	last,
alternativt	alternatively,alternative,
analytiska	analytical,
alternativa	alternative,
tropisk	tropical,
sektion	section,
kubas	cuba,
administrativt	administrative,
monarkin	monarchy,the monarchy,
dömd	sentenced,
administrativa	administration,administrative,administative,
åtal	prosecution,
bin	bin,
dubbelt	double,
bil	car,
teknik	technic,
big	big,
kejsaren	emperor,the emperor,
avlidna	diseased,deceased,
af	of,
möttes	met,
bit	piece,
indonesiska	indonesian,
planeterna	planets,the planets,
rené	rene,
grå	gray,grey,
kolonialtiden	the colonial times,colonial period,
princip	principle,principal,
möjlig	possible,
brett	broad,
stränga	severe,
kristina	kristina,
tillstånd	state,to the dental,condition,
figurerna	figures,characters,
google	google,
identisk	identical,
egyptiska	egyptian,
tolkningar	interpretations,
back	reverse,
historisk	historical,
studerar	study,studies,
cocacola	coca cola,coca-cola,
lars	lars,
västergötland	västergötland,
flygplatser	airports,
måste	have to,must,
lasse	lasse,
per	per,
pratar	talks,talking,
självstyre	autonomy,self-governance,self-government,
saab	saab,
lösningen	the solution,solution,
därför	because,therefore,
nordamerika	north america,
resande	travelers,travelling,
vasaloppet	vasaloppet,
påven	the pope,pope,
ockuperade	occupied,
britannica	britannica,
korta	short,
värmestrålningen	heat radiation,
fallit	fallen,fall,
jimmy	jimmy,
grammy	grammy,
styrelse	board,board of directors,
barcelonas	barcelona,
steven	steven,
brita	brita,
ontario	ontario,
framträdde	emerged,
ökningen	increase,
dalar	valleys,
turkiska	turkey,turkish,
medvetande	consciousness,
jaga	course,hunt,
serie	series,cartoon,
konsul	consul,
bostäder	residences,housing,
torsten	torsten,
jonathan	jonathan,
skillnaden	the difference,
ledningen	conduit,the lead,
mångfald	diversity,variety,
planet	planet,
smycken	jewlery,
sultanen	sultan,
planer	plans,
amfetamin	amphetamine,
skillnader	differences,
reggaen	reggae,
jordbävningen	earthquake,
reidar	reidar,
titel	title,
expedition	caretaker,expidition,expedition,
förbjudna	forbidden,prohibited,
hjärnans	brain,
tropiskt	tropical,
tropiska	tropical,
materia	matter,materia,
tyskland	germany,
eller	or,
voltaire	voltaire,
familjer	families,
årstiderna	seasons,the seasons,
familjen	the family,family,
betalar	paying,
makedonien	macedonia,
anser	view,
anses	be,
konspirationsteorier	conspiracy theories,
lena	lena,
utvecklade	oral,
länders	countries',countries,
samla	collecting,collect,
mutationer	mutations,
nådde	reached,
ritualer	rituals,
storkors	the grand cross,
talades	spoken,spoke,
regionala	regional,
sambandet	the connection,connection,
dramatiker	playwright,dramatist,
judisk	jewish,
sorg	grief,
regionalt	regional,regionally,
agnes	agnes,
uppgår	is,
jason	jason,
stänga	close,off,
stred	fought,
uran	uranium,
frankrike	france,
förut	requires,
sigmund	sigmund,
övergav	abandoned,
intensivt	intensive,hard,
privat	private,
lilla	small,
tillämpningar	applications,
landslaget	the national team,team,
betrakta	view,
sydafrikanska	south african,african,
sahlin	sahlin,
konsten	art,the art,
intensiva	intensive,
kollaps	collapse,
atlas	atlas,
graven	the grave,grave,
passiv	passive,
luleå	luleå,
plikt	duty,
släppte	released,
tjänade	earned,
varnade	warned,
färöarna	the faroe islands,
nonsporting	non sporting,
svts	svts,
tävlingar	competitions,contests,
exemplet	the example,example,
knight	knight,
joel	joel,
ände	end,
slutade	quit,ending,
madeira	madeira,
warszawa	warsaw,
naturens	nature's,nature,
joey	joey,
förlust	loss,
störtades	overthrown,
överhöghet	supremacy,
utbredda	widespread,spread,
vanligaste	frequent,
påsken	easter,
höjdpunkt	climax,high point,
carlo	carlo,
sträcker	stretches,extend,
går	is,goes,
chicago	chicago,
spåras	trace,
tillkomst	origin,established,advent,
senare	later,
sauron	sauron,
placering	position,placement,
börje	börje,borje,
analsex	anal sex,
och	and,
öar	islets,
extremt	extremely,
börja	start,
extrema	extreme,
isländska	icelandic,
mottagaren	the recipient,receiver,
populäraste	rated,most popular,
störning	noise,
honom	his,him,
svårigheter	difficulties,
medeltid	medieval,
turkar	turks,
alaska	alaska,
lagts	added,
katolicismen	catholisism,catholicism,
lagförslag	bill,
miljard	billion,one billion,
färgade	colored,
existens	existence,
protokoll	protocol,
uppnår	achieve,reaches,
uppnås	obtained,is achieved,
talare	speakers,spoke,
privata	private,
stundom	sometimes,somtimes,
når	reaches,
nås	reached,is reached,
filippinerna	filipinos,the philippines,
betraktas	considered,
betraktar	regard,sees,
ovan	above,
lima	lima,
somrarna	the summers,summers,
skivbolag	record company,
kinesisk	chinese,
skotsk	scottish,
chi	chi,
gruppspelet	group stage,group play,
fånga	capture,capturing,
nobel	nobel,
döpt	baptized,
söder	south,
geografisk	geographic,geographical,spatial,
titanics	titanic's,titanic,
konkurrens	competition,
prinsen	prince,the prince,
ledamöterna	commisioners,
förstå	understand,understandable,
utropade	exclaimed,cried out,
bakterier	bacteria,
självständighet	independence,
avsikten	purpose,
iii	iii,
engels	engels,
ansvaret	responsibility,
britney	britney,
tunnel	tunnel,
gabriel	gabriel,
påbörjas	start,starts,
halt	content,stop,
baserad	based,
kedja	chain,
baseras	based,based on,
baserar	base,based,
baserat	based,
kyrkan	the church,church,
väldet	the rule,
fotosyntesen	photosynthesis,
titlar	titles,
do	do,
mozarts	mozart's,mozart,
förlängning	extension,
cecilia	cecilia,
fett	fat,
democracy	democracy,
internationellt	international,internationally,
lanserade	introduced,launched,
internationella	international,
tjänst	service,
vilhelm	vilhelm,
revs	described,
böckerna	books,
rousseau	rousseau,
riktig	real,
klar	clear,done,
billiga	cheap,
föddes	was born,
herrlandskamper	herrlandskamper,men's international contest,
mötte	motte,met,
spannmål	grain,
förbundskapten	manager,
klan	clan,
gammal	old,
terrier	terrier,
finländska	finnish,
rådhus	town hall,courthouse,
förekommit	occurred,
grannar	neighbors,
registrerade	data,noted,
olyckan	incident,
alltjämt	remains,
omslaget	the cover,
halvklotet	hemisphere,
strid	conflict,
matematiken	mathematics,
georg	georgian,georg,
innebär	means,
industrier	industries,
le	le,
la	la,
variationer	variations,
bryts	breaks,
föreställer	depicts,
weber	weber,
dag	day,
avsedda	intended,
spektrum	spectra,
utfärdade	issued,
dam	dam,
dan	dan,
valet	selection,the election,
avslöjar	reveals,
tillkommit	been,accured,
periodiska	periodic,
das	das,
sammanhanget	context,
tolkade	interpreted,
day	day,
kontinuerligt	continuous,continous,
beslut	decision,
morris	morris,
newtons	newton,newton's,
syftade	alluded to,aiming,
emo	emo,
lysande	brilliant,illuminating,
engelskspråkiga	english-speaking,
juridisk	legal,
krita	chalk,
humanism	humanistic,humanism,
pitts	pitts,
kristiansson	kristiansen,kristiansson,
dokumentär	documentary,
inspirerade	inspired,
segern	victory,
programmet	program,the application,
arbetskraft	workforce,labor,
fattigdomen	poverty,
nödvändiga	essential,
matt	dull,
mats	mat's,attention,
kärnan	core,
ren	clean,
deras	their,
försäkra	make sure,
red	eds,
återta	retake,regain,
filmatiseringen	film version,
roterande	rotating,
frank	franks,
webbplats	website,site,
franz	franz,
odlas	cultured,
arbetare	workers,
ronald	ronald,
längre	longer,
inleds	starts,start,
fart	off,speed,
efterträddes	succeeded,
medelhavsområdet	the mediterranean region,the mediterranean area,
referenser	references,
farbror	uncle,
fotografier	photographs,
nivå	level,
south	south,
liberaler	liberals,
stämmer	correct,
genomgår	undergoes,
pga	due,
uppges	reported,
uppger	states,state,
innehålla	include,
insikt	recognition,
därav	thereof,
fruktade	feared,
omständigheter	event,circumstances,
veckan	the week,
leder	leads,
utlopp	outflow,outlet,
energikällor	sources of energy,
kantonerna	cantons,
förklara	explain,declaring,
maidens	maidens,
leden	hinge,lines,the route,
palestina	palestine,
demonstrationer	demonstrations,
bundna	tied,bonded,
släktet	the genus,
stället	instead,the place,
ställer	set,
innehade	held,possessed,
firades	celebrated,was celebrated,
pågående	current,
sjögren	sjögren,
ledamöter	commissioners,
släkten	genera,the family,
ställen	places,
bevarats	protected,preserved,
beskrivningen	description,
domaren	judge,the judge,
matematisk	mathematical,mathematic,
uteslutande	exclusivly,only,exclusively,
kvalificerade	qualifying,
universum	universe,
mälaren	mälaren,
premiär	prime,premiere,
havs	sea,
aristoteles	aristoteles,aristotle,
biologiska	biological,
följd	following,
älgar	moose,
följa	follow,
basist	bassist,
uganda	uganda,
idag	today,
rådande	prevalent,
följt	followed,
följs	followed,
låt	let,
mil	swedish miles,
min	my,
mia	mia,
fötter	feet,on its feet,
kroppar	bodies,
tidningar	press,magazines,
mig	me,
mix	mix,
låg	low,
experter	experts,
besättningen	crew,
lån	loan,
konstverk	work of art,artworks,
konkurrerande	competing,
resurser	resources,
resultatet	the result,result,
dinosaurier	dinosaurs,
varandras	each others,each other,
missionärer	missioners,missionaries,
resultaten	the results,results,
sedan	since,
sist	finally,last,
herman	herman,
liknade	looked like,similar,
stranden	shore,
upprustning	renovation,
irakkriget	iraq war,
republikanska	republican,
rörelsens	movements,movement,
milano	milano,
deuterium	deuterium,
tidskrift	newspaper,magazine,
definiera	defining,define,
viktigaste	most important,
styrka	power,
utgångspunkt	starting point,point of departure,
högtider	holiday,
text	text,
charles	charles,
inhemsk	domestic,native,
ugglas	owl,ugglas,
fungerade	thought,working,
kurfursten	elector,
rumänska	romanian,
järnvägen	railroad,rail,
euroområdet	eurozone,euro area,
rytmiska	rhythmic,
satan	satan,
shahen	the shah,shah,
säker	safety,
bryssel	brussels,
organiska	organic,
snitt	on average,average,
arean	the area,area,
förändrades	changed,
buddhismen	buddhism,buddism,
överlägset	far,
förstår	understand,
regimen	regime,
uppehåll	residence,hiatus,
richards	richards,
idéerna	ideas,
vinsten	the win,gain,
organ	body,
županija	country,
nazitysklands	nazi germany's,nazi germany,
vinster	gains,
majoriteten	the majority,
lyckade	successful,
byggdes	was,was built,
ronaldo	ronaldo,
militärer	military,
krävdes	were required,
national	national,
svenska	swedish,
kapitalet	capital,
svenskt	swedish,
först	first,
egentlig	actual,
debutalbumet	the debut-album,debut album,
reform	reform,
redan	has already,
konverterade	converted,
intog	seized,occupied,took,
carlsson	carlsson,
wembley	wembley,
bör	should,
terräng	terrain,off,
ordentligt	properly,firmly,
översikt	overview,
koncept	concept,
industrialisering	industrialization,
uppskattade	estimated,appreciated,
listan	the list,
hårdare	harder,tougher,
säkerheten	the security,safety,
översättas	translated,be translated,
viktigare	important,more important,
läsning	read,
hämtade	taken,brought,
buddhas	buddha's,buddhas,
empathy	empathy,
miniatyr|karta	thumbnail map,miniature|map,
återförening	reunion,
litteratur	literature,
aktuellt	relevant,
kommunicerar	communicates,
kröntes	crowned,
aktuella	current,
kommendör	commandor,commander,
sachsen	saxony,
fester	celebrations,parties,
inneburit	meant,
befogenhet	warrant,authority,
utsågs	was,was appointed,
medicinsk	medical,
elektroner	electron,
news	news,
ad	ad,
västmakterna	western powers,
tunisien	tunisia,
grupperingar	groups,grouping,
slippa	avoid,
gaza	gaza,
igen	recognize,back,
asteroider	astroids,asteroids,
genomsnittlig	average,
stationen	station,
stationer	stations,
orange	orange,
deep	deep,
thåström	thåström,thastrom,
an	an,
augusti	august,
bruket	use,the use,
stalin	stalin,
ar	is,
ocheller	and/or,
betraktade	watched,
externa	external,
kväve	nitrogen,
tagits	taken,
flyktingar	refugees,
betalade	payed,paid,
fördrag	agreement,treaty,
partner	partner,
prosa	prose,
utom	out,
händelserna	the events,events,the happenings,
lämnade	did,left,
wolfgang	wolfgang,
blodtrycket	the blood pressure,blood pressure,
sångerna	song are,the songs,
omedelbart	immediately,immediate,
heinrich	heinrich,
hinduismen	hinduism,
kallad	called,
kontrollera	control,controlling,
framförallt	above all,
helsingborgs	helsing borg,
kallas	called,
kallar	call,calls,
center	center,
öde	fate,
seth	seth,
antonio	antonio,
sett	seen,
hoppas	hope,
omgångar	cycles,
undvika	avoid,
position	position,
deltar	part,participates,
stores	great,the great's,
kontaktade	contacted,
passade	suiting,suited,
mystiska	mysterious,mystical,
wagner	wagner,
misshandel	assault,abuse,
dagar	day,days,
flertal	majority group,
bevarade	preserved,
vanligt	usual,normal,
hamburg	hamburger,
kampf	kampf,
reformer	reformers,reforms,
lake	lake,
mentala	mental,
landområden	land areas,
streck	bar,
belgrad	belgrade,
förnuft	reason,
uppmärksamhet	attention,attantion,
uppträder	occur,performs,
dubai	dubai,
koden	the code,code,
innehöll	containing,
tusentals	thousands,
likt	like,
journalist	journalist,
works	works,
uppträda	occur,
gudomlig	divine,
albumets	album,album's,
starkaste	the strongest,
värt	worth,
etablerades	established,was established,
minsta	minimum,
est	est,
joachim	joachim,
katarina	katarina,
löser	solve,
skildrar	depicts,
skildras	is depicted,depicted,
gisslan	hostages,
internationalen	international,
definitionen	the definition,
nattetid	overnight,
definitioner	definitions,
starkare	strong,stronger,
leopold	leopold,
arterna	the species,species,
about	about,
socker	sugar,
ärkebiskopen	archbishop,
glada	happy,
mäktigaste	powerful,
tomt	empty,blank,
andel	percentage,share,
anden	spirit,
folkräkningen	census,
medverkar	contributes,contribute,
alexanders	alexanders,
förstärka	strengthen,enhance,
socken	parish,
omgiven	surrounded,
potatis	potato,
monarken	the monarch,
världsliga	worldly,
ljusare	lighter,
föredrar	preferred,
vimmerby	vimmerby,
hatar	hate,hates,
densamma	the same,same,
skog	wood,
kuben	cube,the cube,
strävhårig	hispid,wirehaired,
föga	little,
flyg	flight,airforce,
kärnor	core,
kväll	evening,
klockan	clock,o'clock,
civilbefolkningen	the civilian population,
ryssarna	russians,
brand	fire,
bröder	brothers,
ersättning	replacement,
flygvapnet	air force,
kraft	power,
bud	bid,bids,
vetenskap	science,
utrymme	space,
arbetsgivaren	employer,
lissabon	lisbon,
australiens	australia,australia's,
nedre	lower,bottom,
innanför	inside,
minuter	minutes,
bytet	the exchange,change,
hästens	horses,horse,
circus	circus,
paraguay	paraguay,
tolkningen	interpretetation,interpretation,
omloppsbanor	orbits,
autism	autism,
betydande	important,significant,
vinner	gaining,wins,win,
manlig	male,
särskilda	special,
proteinet	the protein,
proteiner	proteins,
uppfattar	percieves,
picchu	picchu,
stimulans	stimulation,stimulating,
betonade	emphasized,
endast	merely,only,
försämrades	decreased,worsening,
uppfatta	perceived,perceive,
sjön	lake,
tämligen	rather,fairly,
astronomi	astronomy,
variation	diversity,variety,
koncentrationsläger	concentration,concentration camp,
akademisk	academical,
ärkebiskop	archbishop,
cirkel	circular,
philips	philips,
fakta	fact,
winnerbäck	winnerback,
baker	baker,
svag	weak,
uppfattningen	comprehension,view,
framför	in front of,particularly,
förbundet	the union,association,
okänd	unknown,
mäktiga	powerful,
brottslingar	criminals,
slogs	fought,was,
båt	boat,
resor	travels,travel,
påsk	easter,
arkitekt	architect,
antisemitiska	antisemetic,antisemitic,
ozzy	ozzy,
granskning	review,
anfallet	the attack,attack,
upphör	end,
paris	paris,
tillväxten	growth,
deltagit	part,participated,
kapacitet	capacity,
under	for,under,
läge	mode,
svårare	difficult,
nordost	the northeast,
pommern	pommern,
ägande	owning,
jack	jack,
ovanstående	above,
tagit	taken,
utmärks	characterized,
utmärkt	excellent,
öppna	open,
plural	plural,
venus	venus,
matematik	mathematic,mathematics,
verklig	real,
reklam	advertising,advertisement,
parten	party,
markerar	selects,
kropp	body,
bönderna	farmers,
manus	script,
läget	location,
indierna	indians,
läger	camp,
stridigheter	oppositions,strife,
aktivt	active,
drivande	drive,driving,
ebba	ebba,
notera	note,
liberty	liberty,
aktiva	active,
sund	healthy,sane,
kub	cube,
disney	disney,
egyptens	egypt,
språken	languages,
prata	talk,
flera	multiple,
medelhavsklimat	mediterranean climate,
utredning	investigation,
beck	beck,pitch,
parlamentariska	parliamentary,
preparat	substance,
studio	studio,
rysk	russian,
sommartid	summer-time,summer,during summer,
komplex	complex,komplex,
forum	forum,
lagras	stored,
ty	for,
precis	precisely,just,
proportioner	proportions,
svante	svante,
gällande	current,regarding,
koloniserades	is colonized,colonized,
upptäckter	discoveries,discovery,
upptäcktes	discovered,
julie	julie,
erektion	erection,
julia	julia,
övers	transl,
nazistiska	nazi,
misslyckats	failed,
upptäckten	discovery,
försvarsmakt	armed forces,
eftervärlden	the world,
volym	volume,
mattias	mattias,
klassas	classified,
vinst	profit,win,
miniatyr|px|en	miniature,
konserterna	the concerts,concerts,
skicka	send,
behandlingar	treatments,
romaner	novels,
återstående	remaining,
muse	muse,
övertala	convince,persuade,
ludvig	ludvig,
ansökte	applied,
världsarv	world heritage,
fermentering	fermentation,
rörelse	movement,
belgiens	belgium,
igelkottens	the hedgehog's,hedgehog,
henri	henri - it's a name,henri,
mm	millimeter,
arméns	the army's,arm,
antiken	the ancient world,antiquity,
mr	mr,
johanssons	johansson,
utgick	started,
partiets	the party's,parties,
ghana	ghana,
sträckan	distance,the distance,
utlöste	triggered,
trädgård	garden,
florida	florida,
genomfördes	was,was carried out,
fröken	miss,
ena	one,
end	end,
smält	melted,
undantag	except,
väpnade	armed,
ens	even,
gata	street,
elektriskt	electric,
elizabeth	elizabeth,
beskrev	depicted,described,
målen	cases,goals,
förståelse	understanding,
mest	most,mostly,
västvärlden	west,western world,
målet	target,the target,
miniatyr|px|ett	miniature,
elektriska	electrical,
frågade	asked,
 cm	centimeters,cm,
nagasaki	nagasaki,
kategorier	categories,
kubanska	cuban,
beteenden	behavior,
kontrollen	control,the control,
existera	exist,
beskrivit	described,
arbetar	work,works,
kejsare	emperor,
kampen	the fight,fight,
over	over,
arresterades	was arrested,
vitt	white,widely,
besittningar	holdings,possessions,
synonymt	synonymously,
frivillig	optional,
vita	white,
expansion	expansion,
bibelns	the bibel's,
brinner	on fire,
edith	edith,
nytt	new,
dött	dead,
blott	merely,only,
dem	those,
senast	last,
produktion	production,
upptagen	busy,occupied,
livstid	life span,
ansvarar	charge,
jämförelser	comparison,
detroit	detroit,
ersattes	was replaced by,
ställdes	prepared,
newport	newport,
storlek	size,
ursprungligen	initially,originally,
växter	plants,
önskemål	requests,demands,
gymnasium	high school,
group	group,
dessförinnan	before,
träffade	met,
innehållande	containing,
platina	platinum,
nio	nine,
behövs	required,is needed,
kuwait	kuwait,
receptorer	receptors,
användningen	use,the use,
ammoniak	ammonia,
hemland	homeland,
riktning	direction,
danmarks	denmarks,denmark's,
paulus	paulus,paul,
got	got,
stödja	support,
independence	independence,
smala	narrow,
snuset	snuff,
icke	non,
värnplikt	military service,
kandidat	candidate,
fred	peace,
statsöverhuvud	head of state,
undervisade	taught,
samlade	collected,
inom	within,in,
drygt	good,approximately,
statsministern	prime minister,head of state,
studera	study,
tolerans	tolerance,
bredvid	beside,next to,
vetenskapliga	scientific,
samhälle	society,
befolkade	populated,
vetenskapligt	scientifically,scientific,
transporterar	carrying,transports,
transporteras	is transported,
nyheter	news,
säsong	season,
museet	the museum,museum,
museer	museums,musser,
föreslagits	suggested,was suggested,
nhl	nhl,
institutioner	institutions,
rikaste	the richest,richest,
tillåts	is allowed,allowed,
yngsta	youngest,
sexuella	sexual,
nyheten	news,
mercury	mercury,
vikingar	vikings,
tor	thu,
yngste	youngest,
punkten	point,
merkurius	mercury,
å	on,
konventioner	conventions,
ton	tonne,tone,
punkter	points,seq,
tom	tom,
uppkommit	generated,arisen,
tog	was,took,
fördes	out,
adjektiv	adjective,
ifrågasatts	is questioned,questioned,
livealbum	live album,
skildes	separated,was seperated,
meddelande	message,
rädsla	fear,
fördel	advantage,
kulturarv	cultural heritage,
territoriella	territorial,
slutsats	conclusion,
mjölk	milk,
uppmuntrade	encouragement,encouraged,
bridge	bridge,
rad	line,range,
nedgång	decline,decreases,fall,
tänka	thinking,think,
rak	straight,
somliga	some,
störningar	disorder,
växer	growing,grows,
ras	race,ras,
adhd	adhd,
tycks	appears,
tänkt	expected,
industriellt	industrially,industrial,
hittats	found,
kvällen	the evening,
situationer	situations,
lanseringen	the release,
användning	use,
öarna	the islands,
industriella	industrial,
academy	academy,
situationen	situation,
mekaniska	mechanical,
grundskolan	elementary school,
tvingas	forced,system,
skepp	vessel,
elektricitet	electricity,
fralagen	the fra law,
motsatt	opposite,
tanzania	tanzania,
metal	metal,
sekt	sect,
metan	methane,
sjöar	lakes,parks,
inflytande	influence,
flod	river,
utkanten	the outskirts,
dyrare	more expensive,expensive,
idrott	sport,sports,
saga	saga,
järnvägarna	the railways,railways,
queen	drottning,
gränserna	borders,limits,
radio	radio,
earth	earth,
sagt	said,
radie	radius,
absolut	absolute,
skada	damage,
claude	claude,
florens	florence,florens,
vinna	win,
institution	institution,
ägare	owner,owners,
gods	domain,
holländska	dutch,
publik	audience,public,
återstår	remains,
andras	others,
representerade	represented,represent,
mängd	amount,laden,
kommunisterna	communists,the communists,
guatemala	guatemala,
franska	french,
gogh	gogh,
haiti	haiti,
sträckor	distances,
ålder	age,
taubes	taubes,
ändras	be changed,change,
ändrar	change,
ursäkt	excuse,
ändrat	changed,modified,
lovat	promised,
publicerades	published,
tidningen	the newspaper,journal,
utvisning	penalty,expulsion,
kroppen	body,the body,
sakta	slowly,
ockuperat	occupied,
fördomar	bias,prejudices,
kristendomen	chritianity,christianity,
utformade	formed,
behålla	container,
mur	wall,
antikens	ancient,
populär	popular,
slottet	castle,the castle,
finger	finder,
förstås	course,
allra	most,
mun	mouth,oral,
herding	herding,
förhållande	in relation,ratio,
ordnade	arranged,parent,
betonar	emphasize,
omvänt	vice versa,
maniska	manic,
seden	the seed,custom,
dödsorsaken	cause of death,
bildriksdagsval	image election,
nummer	number,
store	great,
kreativitet	creativity,
autonomi	autonomy,
verka	operate,appear,
lösningsmedel	solvent,
läggs	is,
farliga	dangerous,
allierades	allied's,allied,
begränsade	restricted,
förbränning	combustion,
viruset	virus,
lägga	put,add,
november	november,
hitler	hitler,
solljus	sun light,sunlight,
skapades	generated,
rumänien	romania,
reglera	controlling,expell,
möjliggjorde	made possible,allowed,
hastighet	speed,
diktatorn	the dictator,dictator,
homosexuell	homosexual,
skalan	scale,
öster	east,
modernare	mor modern,more modern,
anspråk	claim,
spritt	spread,
drömmar	dreams,
invasionen	invasion,the invasion,
älgen	moose,
n	n,
petrus	petrus,
schizofreni	schizophrenia,
depp	depp,
förståelsen	the understanding,
claes	claes,
della	della,
nationer	nations,
viking	viking,
spelades	filmed,
darwins	darwin,
därigenom	by which,thus,thereby,
vojvodskap	voivodships,voivodeship,
brott	crimes,
anlände	arrived,
känsliga	susceptible,1st&2nd: fragile 3rd: sensitive,
nationen	the nation,
kartan	the map,map,
vanföreställningar	delusions,
varefter	whereafter,
väljs	selected,
ernman	ernman,
äger	owns,
erhållit	obtained,
ökade	increased,
ersatte	substituting,
pekat	pointed,identified,
negativ	negative,
welsh	welsh,
hundra	one hundred,
formatet	the format,size,
ersatts	replaced,
återvände	returned,returning,
återvända	return,
gudom	deity,
dylan	dylan,
generna	the genes,
charlie	charlie,
spelad	played,
tillkännagav	announced,
svavel	sulfur,
kemikalier	chemicals,
fattigare	poorer,
louisiana	louisiana,
jean	jean,
spelat	played,
spelas	played,
spelar	gaming,
mytologin	mythology,
kraftigt	heavily,
järn	iron,
ämnen	agents,
torah	torah,
graden	rate,
europaparlamentet	the european parliament,european parliament,
grader	degrees,
engelskans	english,
utföras	be,performed,
kolväten	hydrocarbons,the hydrocarbon,
kalifornien	california,
använt	using,used,
värnpliktiga	conscripted,inductees,
gavs	was,
belagt	coated,
eld	fire,
grundaren	the founder,founder,
aktiv	active,
regionerna	regions,
ekonomin	the economy,economy,
 au	au,
benämning	term,name,title,
donau	danube,
ämnet	substance,subject,
tillgänglig	available,provided,
protesterade	protested,
auktoritet	authority,
omvärlden	world,surrounding world,
gift	married,
såväl	both,
ladda	load,
modersmål	native language,
bosnienhercegovina	bosnia-hercegovina,
specifik	specific,
tillåtna	allowed,
fotbollen	soccer,
hund	dog,
gifter	marries,
lagstiftningen	law-making,legislation,
enat	united,
hanhon	he/she,male-female,
hushåll	household,
besöka	visit,
jennifer	jennifer,
malaysia	malaysia,
donald	donald,
besökt	visited,
saturnus	saturn,
skapa	create,creating,
estetik	aesthetics,
ultraviolett	ultraviolet,
totalt	complete,wholly,
användare	users,
gösta	gosta,
icd	icd,
diktatur	dictator,dictatorship,
utse	appoint,name,
totala	total,
karaktäriseras	characterizes,is characterised,
elitserien	elite series,elitserien,
monoteism	monotheism,
ishockeyspelare	ice hockey player,hockey players,
tillbringar	spends,
män	males,men,
spelare	player,
hotellet	the hotel,hotel,
meyer	meyer,
titeln	the title,
tvingades	forced,had,
systrar	sisters,
omgången	round,
plus	plus,
internationell	international,
tydliga	clear,obvious,
genomslag	impact,breakthrough,
primitiva	primitive,
civil	civil,civilian,
menade	meant,said,
systemet	the system,system,
tydligt	clear,obvious,
isberg	ice berg,iceberg,
sinne	mind,
anorexia	anorexia,
oförmåga	inability,failure,
omges	surrounded,
omger	surrounding the,
lagt	laid,added,
kjell	kjell,
sicilien	sicily,
gia	gia,
metabolism	metabolism,
wittenberg	wittenberg,
dialekterna	dialects,
fadern	the father,
skulden	the guilt,
barrett	barett,
fängelsestraff	imprisonment,prison,
italien	italy,
skulder	debts,debt,
finns	there is,
eventuell	any,
fusionen	merger,
amerikanerna	americans,the americans,
värvade	recruited,referred,
tillika	also,well,
araber	arabs,
regler	rules,
trio	trio,
bildt	bildt,
hamn	harbor,port,
tronen	throne,the throne,
kambodja	cambodians,
förbud	ban,prohibiting,
liberalism	liberalism,
tätorten	conurbation,agglomeration,
ni	you,
margareta	margareta,
no	no.,
tillverkade	manufactured,
when	when,
nf	nf,
finna	found,
ny	new,
tio	ten,
lösas	solved,
nr	number,no,
tätorter	conurbation,
nu	now,
picture	picture,
phoenix	phoenix,
sätts	is,is placed,
miscellaneous	miscellaneous,
gäster	guests,
tunna	thin,
sätta	insert,
kronprins	crown prince,
väckte	awakened,aroused,
beroendeframkallande	addictive,
vietnam	vietnam,
rom	rome,rom,
ron	ron,
rob	rob,
rod	rod,
dvärg	dwarf,
roy	roy,
koreanska	korean,
udda	odd,
fiktiv	fictitious,
laura	laura,
mottagarens	the reciever,the receivers,
konstitutionell	constitutional,
bär	carryng,berries,here,
tanke	light,in light of,
federation	federation,
även	also,
varvid	in which,
underhållning	entertainment,
flytt	escaped,fled,
krossa	crush,crushing,
metod	method,
inlärning	learning,
hawaii	hawaii,
christmas	christmas,
olyckor	accidents,
lever	liver,
tillverkningen	production,the production,
försvara	defending,
införandet	introduction,the introduction,
trend	trend,
stilar	styles,
kategorirock	category:rock,
colin	colin,
svartån	svartån,
förorter	suburbs,
port	gate,port,
uppgifterna	data,
ifråga	with regards to,challenged,
passa	match,
ögat	eye,
cykel	bicycle,cycle,
månaderna	months,
angelina	angelina,
gräs	grass,
gravitation	gravitation,gravity,
kamp	struggle,fight,
vindkraftverk	wind turbine,
enkla	simple,single,
metaller	metals,
eiffeltornet	the eiffel tower,
turister	tourists,
dublin	dublin,
sina	their,his,
lokal	local,
ankomst	arrival,
asterix	asterix,
tilltagande	increasing,
rafael	rafael,
luften	air,
sikt	term,
etablera	establish,up,
modellen	the model,
trummor	drums,
bolaget	company,the company,
ungerska	hungarian,
russell	russell,
ande	of,spirit,
samfundet	association,
lp	lp,
anda	spirit,
inblandade	involved,
andy	andy,
kurder	kurds,
australian	australian,
turné	tour,
crüe	crüe,
veckorna	weeks,
typerna	the types,
cant	cant,
staten	state,
kär	in love,
övergå	transition,transend,
palestinsk	palestinian,
årets	year,
efterhand	post,
piano	piano,
styras	steered,
drabbades	affected,where hit by,
julius	julius,
musikaliska	musical,
rådgivare	counsellor,advisor,
valla	valla,wax,
jude	jew,
allvarlig	serious,
judy	judy,
humle	hops,
generell	general,
karibiska	caribbean,
musikaliskt	musical,musically,
anpassat	adapted,
uppväxt	growing up,
bönorna	bean,beans,
dokumenterade	documented,
utdelades	distributed,awarded,
hemligt	secret,
annorlunda	otherwise,
hemliga	secret,
främja	further,promote,promoting,
frivilligt	voluntarily,voluntary,
speglar	mirror,
avrättning	execution,
frivilliga	volunteers,optional,
kina	china,
stöter	thrust,run,
simning	swimming,
regeln	rule,
muslimerna	the muslims,
inriktad	oriented,intent,
etablerat	established,
tvserien	the tv show,television program,
levt	survived,
fascism	fascism,
sydliga	southern,
familjens	the familys,family,
flög	fly,flew,
fenomen	phenomenon,
leva	live,
utrikespolitiska	foreign policy,
väntan	awaiting,waiting,wait,
marknad	market,
beror	is,
stridande	conflict,
representation	representation,
väntas	expected,
faser	phases,
orter	varieties,locations,
kartor	maps,
orten	resort,the suburb,
födelse	date,
komplicerat	complex,complicated,
iberiska	iberian,
fasen	phase,
rapport	report,
fartyg	vessel,
böcker	books,
kämpade	fought,
välja	select,
wallace	wallace,
utvecklingen	development,the development,
organisation	organization,
behandlingen	the treatment,the treament,
klassen	the class,
tjänstemän	officals,officials,
marleys	marley's,marley,
passar	suitable,
hergé	herge,
femte	fifth,
märta	märta,
hamilton	hamilton,
tredjedel	a third,third,
hotar	threatens,
term	term,
opera	opera,
snabb	instant,
namn	name,
futharkens	futharkens,the futhark's,
viggo	viggo,
alternativ	alternative,
hotad	threatened,
färger	color,colors,
bildning	education,form,
semifinal	semifinals,semi finals,
förhandlingarna	negotiations,
stående	standing,
amerikansk	american,u.s.,
åsikt	opinion,
tillhörighet	affiliation,
behandlas	treated,
upprepade	repeated,
accepterad	acceptable,
stortorget	stortorget,
årliga	annual,
profil	profile,
accepterar	accepts,accept,
accepterat	accepted,
kent	kent,
variant	variant,variety,
juldagen	christmas day,
zuckerberg	zuckerberg,
etanol	ethanol,
nått	reached,
hjalmar	hjalmar,
gallien	gaul,
soundtrack	soundtrack,
arbetet	work,the work,
händelse	handel,
traditionen	the tradition,tradition,
motion	exercise,
traditioner	traditions,
place	place,
någonsin	ever,
politiken	policy,the politics,
hemsida	homepage,
blood	blood,
origin	origin,
begår	commits,commit,
såldes	sold,
självbiografi	autobiography,
kontrollerade	controlled,
given	given,
nuvarande	current,
vågor	waves,
okända	unknown,
sydafrika	south africa,
cullen	cullen,
bahamas	bahamas,
skjuter	slide,
givet	granted,given,
folkmängden	population,
personlighetsstörningar	personality disorders,
spelats	recorded,been played,played,
webbplatser	websites,
kronprinsessan	crown princess,
användandet	use,
grund	because,
montenegro	montenegro,
alan	alan,
kallade	called,
hur	how,the,cage,
hus	house,a house,
webbplatsen	the website,site,
population	population,
smeknamn	nickname,
nathan	nathan,
begravning	funeral,
marinen	navy,marines,
löfte	promise,
kontroll	control,
framställning	preparation,production,
modeller	models,
bildades	formed,was formed,
hjärtat	the heart,
rena	pure,
mottagare	receiver,
ana	feel,ana,
anc	anc,
kromosomerna	the chromosomes,
maten	the food,
mando	command,
rent	clean,
jordskorpan	earth crust,
världen	world,the world,
avstånd	distance,
förste	the first,first,
första	first,
fysikaliska	physical,
förhållandena	conditions,the conditions,
gustavs	gustavs,gustav,
kust	coastal,coast,
periodvis	periodically,
stjärnornas	stellar,the star's,
knutna	associated,attached,tied,
diskussioner	discussions,discussion,
falla	fall,
fria	free,
invånarna	residents,
täcks	covers,
lisbet	lisbet,
astronomiska	astronomical,
erkänner	admits,recognize,
stövare	hound,
herren	the lord,
tron	faith,
ronaldinho	ronaldinho,
mänskligheten	humanity,
bernadotte	bernadotte,
isolering	isolation,
sjunka	decrease,descend,
tror	believe,
bandets	the bands,band,
gula	yellow,
guld	gold,
flydde	fled,
motivet	the motive,subject,
ovanligt	unusual,
gult	yellow,
iväg	away,off,
ovanliga	unusual,rare,
analys	analysis,
berättelser	stories,
webbkällor	web sources,
larsson	larsson,
grundandet	founding,
tränaren	coach,
jazz	jazz,
administrativ	administrative,administration,
nedåt	down,
väder	weather,
theta	theta,
forsberg	forsberg,
beredd	prepared,
tränade	trained,
dramat	drama,the drama,
umeå	umeå,
joker	joker,
republika	republic,
osäkert	insecure,unclear,uncertain,
förmån	benefit,
minnen	memories,memory,
underlätta	ease,
kraftigare	greater,
inspelningen	recording,
uppdraget	assignment,
tekniskt	technical,
college	college,
stanley	stanley,
minnet	memory,
älg	elk,moose,
freden	the peace,peace,
federal	federal,
skett	done,happened,
önskade	wished,
hämtar	download,is,
återigen	yet again,
intresserad	interested,
hämtat	collected,taken,
konstnären	artists,the artist,artist,
mellan	between,
konstnärer	artists,
bekämpa	fight,
ruiner	ruins,
dödade	killed,
myter	myths,
summa	sum,
sydeuropa	southern europe,
region	region,
ordagrant	literal,verbatim,
spindlar	spiders,
lenins	lenin,lenin's,
introducerades	introduced,
gjorde	did,
gjorda	made,done,
pakistan	pakistan,
utgåvor	editions,issues,
period	period,
pop	pop,
fransk	french,france,
werner	werner,
statens	state,the government's,
utformning	layout,formation,
hävda	claim,asserting,
poe	poe,
skånska	scanian dialect,scanian,
howard	howard,
folken	the peoples,people,
strikta	strict,
förekomsten	existence,presence,
dagarna	the days,day,
musikstil	music,music style,
folket	the people,people,
invaderade	invaded,
anderna	andes,the andes,
sändebud	envoy,
andres	andres,
stadshus	town hall,
andrew	andrew,
kapitulation	surrender,capitulation,
tiger	silent,
övrig	other,
minister	minister,
epok	epoch,
champions	champions,
använder	uses,
gustafsson	gustafsson,
riktade	targeted,
allsvenskan	headlines,
cash	cash,
arnold	arnold,
spreds	spread,
fiende	enemy,
grundlagen	constitution,the constitutional law,
synvinkel	angle,
universums	universe,
pippi	birdie,pippi,
kuriosa	trivia,
knyta	tie,
grönland	greenland,
status	status,
producera	produce,producing,
republikens	republic,
fysiologi	physiology,
protoner	protons,
persons	a person's,persons,
linjerna	the lines,lines,
göring	goring,cleaning,
privilegier	privileges,
vatikanstaten	vatican city,vatican,
relaterade	related,
modet	courage,
medvetna	aware,conscious,
kommunistisk	communistic,communist,
breda	wide,
hårdvara	hardware,
without	without,
nordkoreas	north korea,
medellivslängd	average lifespan,life expectancy,
arkitekten	architect,the architect,
kopplingen	coupling,
fördelas	distribute,distributed,
listorna	menus,the lists,
kommentarer	comments,
förklarades	was explained,explained,
enligt	according to,
kill	kill,
knäppupp	knäppup,knäppupp,
harrison	harrison,
moçambique	mozambique,
leta	search,check,
utvinns	extracted,
starka	strong,
tim	tim,h,
rose	rose,
regent	regent,
rosa	pink,
utbyte	yield,trade,
blod	blood,
lett	resulted,
pendeltåg	commuter,
delstat	land,
guldbollen	golden ball,guldbollen,
ross	ross,
riket	the land,
mesta	most,
porto	postage,
vampyren	the vampire,vampire,
delhi	delhi,
utrikespolitik	foreign policy,foreign affairs,
uppslagsordet	lookup word,
kille	guy,
tid	time,
majoritet	majority,
inflation	inflation,
vampyrer	vampires,
riken	the kingdoms,kingdoms,
kommentar	comment,
afrikas	africas,
talrika	numerous,
mexikanska	mexican,
cooper	cooper,
anföll	attacked,
rammstein	rammstein,
verksamheten	activity,
innebära	mean,
teorin	theory,the theory,
gång	once,time,
passera	pass,
latinet	latin,
alkoholer	alcohols,
verksamheter	operations,businesses,
försvarare	defenders,defender,
tiders	days',
fiktion	fiction,
inspirerades	inspired,
sitta	sit,
stopp	stop,
moon	moon,
härledas	derived,
lärda	scholars,savants,
buddha	buddha,
lärde	learned,
uppbyggnad	construction,
storhetstid	heyday,
liberala	liberal,
football	football,
servrar	servers,
geografi	geography,
genom	through,
tyskt	german,
mandelas	mandelas,mandela's,
tyska	german,
tyske	german,
förbindelser	relations,
on	on,
om	of,if,
edwall	edwall,
spelet	the game,game,
og	og,
of	of,av,
oc	o.c.,oc,
stand	stand,
os	os,
or	or,
befäl	command,
koppling	clutch,connection,
cambridge	cambridge,
ansträngningar	effort,
domstol	court,
burton	burton,
befinna	be,
mental	mental,
medlemsstaternas	member,member state,
valley	valley,
serbien	serbia,
förrän	until,
jul	christmas,
inriktning	direction,orientation,
ingredienser	ingredients,
manuskript	manuscript,
värre	worse,
ämbetsmän	officers,bailies,
chaplin	chaplin,
kvinnornas	womens,women,
taylor	taylor,
felix	felix,
närmast	closest,
fjorton	fourteen,
pengar	money,
ökning	increase,
operation	operation,
köpenhamn	copenhagen,
många	many,
roses	roses,
utgifter	expenditure,expenses,
regissör	director,
babylon	babylon,
visade	showed,
separata	separate,
grupp	group,
sällskapet	society,the company,
symbol	symbol,
erövring	conquest,
missbruk	abuse,
vinnaren	winner,
observatörer	observers,
symtomen	symptoms,ymptoms,
dog	died,
barcelona	barcelona,
calle	calle,
erfarenhet	experience,
visby	visby,
all	any,
ali	ali,
alf	alf,
separat	seperate,separate,
konsekvens	impact,consequence,
stödde	supported,
samhällen	communities,societies,
utomliggande	outlying,
sakrament	sacrament,
antogs	was assumed,
uppdrag	job,missions,
persiska	persian,
funktionerna	functions,the functions,
kapitulerade	surrendered,
röstade	voted,
ögonen	eyes,
gary	gary,
påstående	claim,assumption,
program	application,
cykeln	cycle,
kvar	left,
löper	runs,at,
färgerna	colors,
woman	woman,
litet	small,
oavgjort	tie,draw,
song	song,
far	father,
fas	phase,
fat	barrel,
runtom	throughout,around,
simpsons	simpsons,
fan	fan,
sony	sony,
unionens	the union's,
tjeckiska	czech,
choklad	chocolate,
knutsson	knutsson,
list	cunning,
ingående	input,enter into,
förtryck	opression,
lisa	lisa,
över	over,
iran	iran,
grekland	greece,
ted	ted,
istiden	ice age,the ice age,
tex	for example,e.g.,
design	design,
haag	the hague,
what	what,
enklaste	easiest,
sun	sun,
vaginalt	vaginal,
kinesiska	chinese,
spelning	gig,
mördades	was murdered,
guns	guns,
fäste	bracket,
christian	christian,
dottern	daughter,
upptäcka	discover,
regerade	reigned,
avrättades	was executed,executed,
leeds	leeds,
fjärdedel	quarter,fourth,
upptäckt	discovered,found,discovery,
norden	the nordic countries,north,
nordens	the scandinavian countries',scandinavia,
upptäcks	discoverd,
råder	advises,is,
kommande	upcoming,
soloalbum	solo album,
kärnvapen	nuclear,nuclear weapons,
tillhörde	belonged to,belonging to,
magnitud	magnitude,
arabemiraten	united arab emirates,
nyfödda	newborn,
påföljande	following,subsequent,
uppkomst	origin,
filmerna	films,the movies,
stöd	support,
syfte	purpose,
syfta	aim,refer,
smak	flavoring,
socialdemokraterna	members of the social democracy,social democratic,
anarkism	anarchism,
succé	succession,
kommittén	the committee,
branden	the fire,
förebild	role model,
autonom	independent,autonomic,
bekräftade	confirmed,
genomsnittliga	average,
israel	israel,israeli,
permanenta	permanent,
alltid	always,
akademiens	academy,the academy's,
glas	glass,
hålet	hole,the hole,
floyd	floyd,
glad	happy,
östra	eastern,
naturligt	natural,
legender	legends,
godkänt	approved,pass,
decenniet	decade,
gatorna	the streets,streets,
decennier	decades,
kryddor	spices,
förhåller	relationship,
naturliga	natural,
pony	pony,
duett	duet,
bosatt	resident,lived,
styrs	ruled,
elektrisk	elektirsk,
historiskt	historic,historical,
court	court,
breaking	breakingpoint,breaking,
brittisk	british,
satanism	satanism,
historiska	historical,
härstamning	lineage,origin,descent,
välgörenhet	charity,
rocksångare	rock singers,rock singer,
taget	time,
sven	sven,
tagen	taken,
grundämne	elemental,element,
fötterna	feet,
ångest	anxiety,
fötts	born,borned,
atomer	atoms,
regnar	rains,
anarkistiska	anarchist,
praktiska	practical,
bildade	formed,
tsar	tsar,
homosexuella	homosexual,gay,
grande	grande,grand,
greklands	greek country,
människors	humans,human,
instabil	unstable,
längs	along,
september	september,
sträckte	extended,
emmanuel	emmanuel,
mission	mission,
australien	australia,
längd	length,
retoriska	rhetorical,
islam	islam,
lyder	reads,obeys,
rika	rich,
abbey	abbey,
centralort	central city,centralot,
rikt	target,rich,
prag	prague,
stephen	stephen,
argentina	argentina,
jämte	plus,
fenomenet	the phenomenon,phenomenon,
kategorieuropeiska	european category,
styret	gate,
medborgerliga	civil,
kärna	core,quarks,
postumt	posthumously,
landborgen	the ridge,
marcus	marcus,
försöken	attempts,the tries,
journalisten	journalist,the journalist,
forna	former,
stilen	style,
slidan	vaginal,
journalister	journalists,
försöker	tries,trying,
principer	principals,principles,
kustlinje	coastline,
ringar	rings,
drycken	the drink,
betyg	grades,
brother	brother,
aldrig	never,
mongoliet	mongolia,
stenar	stones,blocks,
ollonet	penis head,glans,the glans,
därvid	therewith,
nepal	nepal,
europas	europe,
hill	hill,
väg	way,
kvinna	woman,
väl	good,
vän	friend,
poliser	police,
ökad	increase,increased,
islamistiska	islamist,
ersatt	replaced,
beräknades	calculated,estimated,
kritiserat	criticized,criticised,
bära	carry,mean,
ökar	increases,
polisen	police,
faller	fall,
fallet	case,the case,
stavningen	the spelling,
konsumtionen	consumption,
fallen	case,cases,
aminosyror	amino acids,
filosofins	philosophy,the philosophy,
heinz	heinz,
colombia	colombia,
pablo	pablo,
bland	including,
blanc	blanc,
story	story,
infört	introduced,
lördagen	the saturday,saturday,
automobile	automobile,
misslyckas	fail,fails,
harris	harris,
stort	large,big,
motiveringen	the motivation,ground,
storm	storm,
kristendomens	christianity's,christianity,
stora	large,big,
ecuador	ecuador,
familjerna	families,
mikael	mikael,
gränser	borders,frontiers,
hotel	hotel,
kongress	congress,
serotonin	serotonin,
framtiden	future,the future,
hotet	threat,
fattigaste	the poorest,
gränsen	limit,border,
besökare	visitors,
siffra	number,figure,
king	king,
illegala	illegal,irregular,
matcherna	the games,
direkt	direct,
nöd	distress,emergency,
pjäsen	piece,
dans	dance,
kategorisommarvärdar	category summer hosts,
guden	god,the god,
stjärnan	the star,
tillåta	allowing,
klubb	club,
anläggningar	plants,facilities,
kusin	cousin,
tilldelas	assigned,
omskärelse	circumcision,
slåss	fight,
divisionen	division,
wilson	wilson,
bedriver	operate,
inriktningar	specializations,
dialekt	dialect,
jämförelsevis	comparative,in comparison,
judas	judas,
judar	jews,
kiss	view,
folkgrupper	communities,ethnic groups,
electric	electic,electric,
dagliga	daily,
park	park,
stjärnans	the stars,
dagligt	daily,
industrialiserade	industrialized,
sånger	songs,
mineral	minerals,mineral,
windows	windows,
influensan	the influenza,
sången	the song,song,
borgmästare	mayor,
statsskick	polity,government,
kosovo	kosovo,
tjugo	twenty,
ursprungliga	original,
kolonialism	colonialism,
tilly	tilly,
månen	the moon,
tills	until the,until,
beräkningar	calculations,
canaria	canaria,
bidrog	contributed,
moses	moses,
hit	to here,here,
hiv	hiv,
stormakterna	great powers,
inklusive	including,
vardera	either,each,
fattiga	poor,
händer	happening,hands,
himmler	himmler,
solsystemet	the solar system,
utvidgade	expanded,
tvkanaler	tv channels,
mediciner	medicines,
knapp	button,bare,
tidszon	timezone,time zone,
vincent	vincent,
norrköping	norrköping,
poäng	score,
virginia	virginia,
utsatt	exposed,
bars	bar,
etiopien	ethiopia,
art	kind,art,
bart	offense,bart,
arv	heritage,
fiske	fishing,
bara	only,
arg	angry,
flyttade	moved,
stjäla	steal,
arm	arm,
barn	child,
pär	pär,
bortsett	except,
planeras	is planned,planned,
överföring	transfer,
uppskatta	appreciate,
inga	not,no,
planerat	planned,
planerad	planned,
korea	koreans,korea,
verksamhet	work,activity,
där	where,in which,
intäkter	revenues,incomes,
herrar	gentlemen,men,
uppkom	arose,
godkändes	approved,
tiderna	the times,time,
balkanhalvön	balkan peninsula,
startades	started,
lyssnar	listens,listen,
lägret	the camp,camp,
klassificeras	classified,
hypotesen	the hypothesis,
lära	get to know,
borta	gone,
vidare	moreover,furthermore,
lärt	learned,
stärktes	strengthened,was strenghten,
belägna	located,disposed,
besegrade	defeated,
östtyskland	east germany,
slott	castle,
hypoteser	hypotheses,hypothesis,
ps	ps,p.s.,
java	java,
göteborg	gothenburg,
personalen	personnel,the staff,
kungafamiljen	the royal family,
johannes	johannes,john,
avslutade	ended,finished,
byxor	pants,
resultat	results,result,
ph	ph,
pi	pi,
chandler	chandler,
flight	flights,flight,
togs	taken,were taken,
publiken	audience,
sydafrikas	south african,south africa's,
rättigheterna	the rights,
gården	farm,
konflikter	conflicts,conflict,
konflikten	conflict,
deltog	participated,
sådan	such,
inspelningar	recordings,
ägs	is owned,owned,
styr	controls,
ris	rice,
rik	rich,
sjöarna	the lakes,lakes,
byggnaderna	building,the buildings,
skeppen	the ships,
fysisk	natural,physical,
demografi	demographics,
tidpunkten	the time,the moment,time,
ideologier	ideologies,
sjunkit	decreased,
förföljelse	persecution,
torbjörn	torbjörn,
spears	spears,
låtit	let,had,
bröllopet	the wedding,wedding,
byar	villages,
skåne	skåne,
uppbyggd	structered,structured,built-up,
författare	author,
berömt	praised,
kokpunkt	boiling point,
finansiera	fund,finance,
italiensk	italian,
sjunga	sing,
edge	edge,
vetenskapen	the science,science,
kyrkans	the church's,church,
alfabet	alphabets,alphabet,
uttalande	statement,
komplett	complete,
konstitution	constitution,
remmer	remmer,
dåtidens	past times,that time,
prince	prince,
bidragande	contributors,
folkräkning	census,
skalv	quake,
minoriteter	minorities,
bostad	lodge,property,
omedelbar	instant,immediate,
försvunnit	disappeared,
skall	is,shall,
minoriteten	minority,
idé	ide,
emigrerade	emigrated,
skala	scale,
färdiga	finished,
synnerhet	specially,particular,
djupare	depth,deeper,
begravdes	buried,
användas	used,
stoppade	stopped,
upplevelse	experience,
exakt	accurately,
våldsamma	violent,
näringsliv	business,
banbrytande	groundbreaking,
sammansättning	composition,
hittades	was found,
hittas	found,
minskning	decline,
landskommun	rural municipality,
norrut	north,
sjöfart	sea voyage,maritime,
kongo	congo,kongo,
lettland	latvia,
trummis	drummer,
krigare	warrior,
flottan	the fleet,navy,
thailand	thailand,
huvudstad	capital,
låtarna	the songs,songs,
ungefär	about,
höjden	height,
föräldrar	parents,
grekerna	greek,greeks,
prov	test,
frälsning	salvation,
fungera	act,
anne	anne,
trinidad	trinidad,
anna	anna,
höjder	altitudes,heights,
turism	tourism,
palmes	palme,plame's,
ställningen	position,
tävlade	competed,
presenteras	presented,
anklagades	accused,
judendom	judaism,jewism,
kostnaderna	the costs,
grundläggande	primary,
påtryckningar	pressures,pressure,
tätt	tight,tightly,
virus	virus,
utropades	proclaimed,was proclaimed,
dialog	dialogue,
täta	close,seal,
socialistisk	socialistic,socialist,
oktoberrevolutionen	october revolution,
genomföras	carried out,
medborgarna	the citizens,citizens,
reglerna	rules,
hållet	cohesive,way,
abbas	abbas,
km²	square kilometre,
laget	the team,stroke,
håller	is,holds,
dricka	drinking,
fast	solid,even though,
jugoslavien	yugoslavia,
bagge	bagge,
bruk	using,use,
laila	laila,
ateister	steister,
delning	pitch,
rasade	collapsed,
regionen	the region,region,
längtan	longing,
sköter	handles,handle,
kritikerna	the critics,
delta	delta,
tidigast	the earliest,
junior	junior,
karolinska	caroline,
anklagelser	allegations,
planeternas	the planets,planets,the planets',
världskrigen	the world wars,world wars,
styrande	rulers,governing,
aktier	share,
homo	homo,gay,
guyana	guyana (name),guyana,
tolka	interpreting,interpret,
handels	commercial,
z	z,
tidens	time's,
svenskspråkiga	swedish speaking,
ägdes	owned,
singlarna	singles,
tidpunkt	date,time,
home	home,
däribland	including,
graham	graham,
uppskattningar	estimates,
rainbow	rainbow,
stadion	stadium,
möten	meetings,
höga	high,
psykoterapi	psychotherapy,
operan	opera,
mötet	the meeting,meeting,
hanen	the cock,male,
urval	selection,
skyddas	protected,
skyddar	protects,
sutra	sutra,
beräknas	calculated,
beräknar	computes,values,
tittarna	the viewers,viewers,
medina	medina,
stadigt	stable,steadily,
konvertera	convert,conversion,
betyder	means,
råkar	happens,happens to,
kaspiska	caspian,
modernismen	modernism,
klubbens	club,
oväntat	unexpected,
underlättar	facilitates,
vice	vice,
europeiska	european,
parallella	parallel,
mesopotamien	mesopotamia,
nasa	nasa,
lagstiftning	law-making,regulation,
europeiskt	european,
nash	nash,
förhandla	negotiating,
psykologi	psychology,
beträffande	on,
kanal	channel,
steve	steve,
jimi	jimi,
låter	let,
moseboken	genesis,
kolonialismen	the colonialism,
simon	simon,
uppmaning	call,exhortation,
fortfarande	still,
romerna	the romani,the romani people,
kazakstan	kazakstan,
generellt	generally,
generella	overall,general,
hinduism	hinduism,
fotnoter	footnotes,
pengarna	the money,money,
varierar	varies,
vapen	weapons,weapon,
kategoritvseriestarter	category television series starts,
varierat	varied,
sjukdomar	disease,
medverkade	participated,
kommitté	committee,
avslutas	close,ends,closing,
avslutat	completed,
tvinga	force,
historikern	historian,
äta	eat,
inleder	start,initiates,
noter	notes,notation,
öron	ear,
läkemedel	medicine,
utanför	outside,
melodier	melodies,
byggd	built,
demokratiska	democratic,
bygga	building,build,
indirekt	indirectly,
skadad	damaged,
åtminstone	at least,
århundradet	century,
influerad	influenced,
anderssons	anderssons,
skadas	damaged,
västlig	western,
konstant	constant,
folk	public,people,
influerat	influenced,
hölls	was held,was,
assisterande	assistant,assisted,
kris	crisis,
skrivna	written,
domkyrka	cathedral,abbey,
krig	war,
dramatiska	dramatic,
bröts	was fractured,
insats	stake,
koloni	colony,
hdmi	hdmi,
producenten	the producer,
turismen	tourism,
diamanter	diamonds,
åtgärder	measures,
filosofi	philosophy,
astrid	astrid,
tvingats	forced,had,
buddhistiska	buddhistic,buddhist,
ukraina	ukraine,
metro	metro,
innehar	holds,
innehas	held,
elektronik	electronics,
springsteens	springsteen's,springsteens,
plattan	plate,
fortsätter	continues,
populärkulturen	popular culture,
översättningar	translations,
tjänar	earns,serves,
zlatan	zlatan,
reda	out,find our,
gemenskap	fellowship,community,
föreställande	depicting,
motor	engine,
juryns	the jury's,jury,
redo	prepared,
varpå	whereupon,
from	from,
bestämmelser	measures,conditions,
usa	usa,
fel	errors,
fem	five,
sevärdheter	attractions,
upplöstes	dissolved,
källorna	source,the sources,
inlandet	inland,the inland,
öppnat	opening,
andliga	spiritual,
penis	penis,
införande	introduction,
hindrade	prevented,
vägrade	refused,
reguljära	regular,
beskriva	describe,
automatiskt	automatic,
tar	takes,
tas	is,is taken,
föreslår	suggests,suggest,
platser	points,places,
crick	cricket,crick,
platsen	place,site,
treenigheten	tinity,the trinity,
tag	while,
tal	speech,
kanadensiska	canadian,
sir	sir,
ondska	evil,
löften	promises,
beyoncé	beyoncé,
six	six,
brian	brian,
sig	to,
undantaget	except,
sin	its,
väpnad	armed,
kostym	costume,
kontroversiellt	controversial,
avsnitten	sections,
oavsett	whether,regardless,
tack	thanks,
religiös	religious,
bertil	bertil,
kategoriwikipediabasartiklar	category wikipedia basartiklar,
kontroversiella	controversial,
eritrea	eritrea,
light	light,
centralorter	centers,
kommunikationer	communications,
öresund	Øresund,
jolie	jolie,jolies,
besegrat	defeated,
mekka	mecca,
blandad	blended,
skapande	building,creative,
företrädare	representatives,
elin	elin,electrical,
elit	elite,
karlstad	karlstad,
blandas	mixes,
spotify	spotify,
stiga	rise,rising,
uppmärksammad	attention,noticed,
befolkning	population,
byn	village,
återvänt	returned,returning,
permanent	permanent,
försvar	defence,defense,
lärjungar	disciple,
uppmärksammat	attention,noticed,
carola	carola,
skede	period,analysis,
cypern	cyprus,
verkligen	real,
washington	washington,
fler	more,
andlig	spiritual,
östtimor	east timor,
satelliter	satellite,
exempelvis	e.g.,
komma	access,
billy	billy,
växande	growing,
konungariket	kingdom,
studios	studios,the studio's,
australiska	australian,
säsonger	seasons,
barnets	child,
byter	changes,exchanges,
kvarteret	quarter,the neighborhood,
säsongen	season,
studion	studio,the studio,
kritik	criticism,critisism,
alger	algae,
förbjuda	ban,prohibiting,
uggla	owl,
minskad	decreased,
hantverkare	craftsman,handy worker,
fiktiva	fictitious,
svar	answer,response,
nobelpristagare	nobel laureates,
minskat	decreased,has decreased,
centralamerika	central america,
minskar	decrease,
förutsättningar	prerequisites,condition,
hörs	heard,
hört	heard,heared,
hjälpt	helped,
vulkanutbrott	vulcano eruption,volcanic eruption,
utmärker	characterized,
höra	know,
hjälpa	helping,
york	york,
studioalbumet	studio album,
philip	philip,
domare	judge,
hörn	corner,
fotbollslandslag	football team,national football team,
gångna	past,
anslutning	connection,
tyst	quiet,silent,
waterloo	waterloo,
barns	child,childrens,children,
via	through,
adrian	adrian,
tvserier	tv shows,
tysk	german,
rudolf	rudolph,rudolf,
ovanpå	top,on top of,
revolutionens	revolution,the revolutions,
isbn	isbn,
brasilien	brazil,
velat	wanted,
nietzsches	nietzsche,nietzsche's,
regenter	monarchs,regents,
skyddade	protected,
nätverk	network,
enkelt	easy,
åtskilliga	several,
fågelhundar	bird dogs,
meddelanden	messages,
omfattning	extent,
misslyckande	failure,
sankta	sankta,saint,
diskutera	discussed,
rösträtt	vote,right to vote,
valde	selected,chose,
valda	chosen,
vingar	wings,
juli	july,
vind	wind,
dödligheten	mortality,
resterande	remainder,remaining,
belgien	belgium,
lutning	closing,incline,
holland	holland,
franske	the french,french,
birgitta	birgitta,
tommy	tommy,
framgång	success,
algeriet	algeria,
franskt	french,
tomma	empty,
tyskarna	germans,the germans,
heydrich	heydrich,
fyrtio	forty,
cohen	cohen - it's a name,cohen,
benny	benny,
avgörs	decided,is determined,
blir	become,is,
farligt	dangerous,
ringen	ring,
gäng	group,thread,
intervju	interview,
storbritannien	uk,
byggas	prevented,build,
uppfann	invented,
lopp	race,
ansåg	thought,found,considered,
besittning	dominion,possess,
kristi	kristi,
betydligt	considerably,
centra	center,
ström	power,
centre	centre,
who	who,
intogs	was captured,
staternas	states,
öken	desert,
planerade	planned,
förbundsrepubliken	the federal republic,federal republic of,
undersökte	investigated,
regeringschef	government,
miljontals	millions,
enbart	only,
judendomen	judaism,
kategoriamerikanska	u.s. category,
moberg	moberg,
uefa	uefa,
blandade	mixed,
funktionella	functional,
debatt	debate,
julafton	chistmas eve,christmas eve,
pastoral	pastoral,
komplicerad	complicated,
dödades	were killed,
filmen	the movie,film,
nilsson	nilsson,
filmer	films,movies,
röster	votes,
beroende	dependent,
hållning	position,
allmänhet	in general,general,
träffa	meet,see,
gränsar	adjacent,
överens	in agreement,
gudar	gods,
linje	line,
presley	presley,
hett	hot,
närstående	relative,kindred,
samtycke	consent,
städer	urban,cities,
begäran	request,
förbinder	connects,undertake,
torka	dry,
respektive	and,respective,
mestadels	mostly,
kvinnorna	the women,
berömd	famous,
nationernas	the nations,nations,
rikare	richer,
motståndare	opponents,opponent,
ansågs	was,seemed,
funktion	function,
upplysning	enlightenment,
praktisk	practical,
sydstaterna	southern states,southern united states,
samhället	the society,society,
vandrar	wanders,migrates,
joe	joe,
swift	swift,
jon	jon,
sångaren	singer,
influenser	influence,influences,
ingemar	ingemar,
påtagligt	substantially,markedly,
kolhydrater	carbohydrates,
april	april,
västerländsk	western,
brons	bronze,
vattnets	water,the water's,the waters,
bronx	the bronx,
förespråkare	spokesman,proponent,
betecknar	represents,denotes,
betecknas	denote,
exakta	exact,
korruption	corruption,
wall	wall,
vittne	witness,
publicerad	published,
walt	walt,
cirka	about,approximately,
utsedd	appointed,
styrkor	strenghts,forces,
publiceras	published,
framträdanden	appearances,
publicerat	published,
utkom	issued,
klara	clear,
dödshjälp	euthanasy,euthanasia,
kopplade	connected,
bbc	bbc,
beskrivning	description,
månar	moons,
klart	clear,done,
månad	month,
strindbergs	strindberg's,strindberg,
naturtillgångar	natural resources,
liverpool	liverpool,
nickel	nickel,
försvaret	the defense,
turneringen	the tournament,
dominera	dominate,
lutherska	lutheran,
försvann	disappeared,
hms	hms,
fortsättningen	the continuation,remain,
neutrala	neutral,
deklarerade	declared,
last	load,
plikter	duties,
present	gift,
godkännande	approval,
bråk	fights,fraction,
problemen	the problems,
officiell	official,authentic,
största	biggest,maximum,largest,
anpassa	adjust,
fördelade	divided,distributed,
nominerades	was nominated,nominated,
wild	wild,
madeleine	madeleine,
folktro	folklore,
explosionen	the explosion,
sagan	story,
vuxit	grown,
gemensamt	single,in common,
bosättare	settlers,
syftar	refers,seek to,
motiv	subjects,motif,
jehovas	jehovas,jehova's,
röra	move,
uppstå	develop,
ramels	ramel's,
halv	half,
buddhism	buddhism,
pojkar	boys,
samband	connection,
inch	inches,
skickade	sent,
gett	gave,
annekterade	annexed,annexation,
tvister	conflicts,disputes,
mottagande	host,
övervägande	predominant,predominantly,
romeo	romeo,
romer	romani people,roma,
student	student,
raka	straight,
rätt	entitled,
misstag	error,mistake,
klubbar	clubs,
vilar	rests,
banden	bands,the bound,
terrorismen	terrorism,the terrorism,
undersökningar	studies,
närma	approach,approximate,
ekosystem	ecosystem,
övertyga	convince,
bandet	band,
organisationens	organization,the organizations,
hårdrocken	hard rock,
lön	salary,
biologisk	biological,
möjligheter	potential,
uppkommer	arises,
möjligheten	the ability,
rachels	rachel's,
erfarenheter	experiences,experience,
högskolor	colleges,
förtroende	confidence,
miljöer	environments,
antisemitism	antisemitism,
rocken	rock,
brutit	broken,
mytologiska	mythological,
jarl	earl,jarl,
genombrottet	breakthrough,
alldeles	completely,altogether,
hoppa	drop out,
bell	bell,
sky	sky,
rättsliga	legal,
engelsk	english,
ske	be,happen,
ska	will,
fyller	turns,
sanskrit	sanskrit,
färgen	color,the color,
olle	olle,
agerande	behavior,
älska	love,
know	know,
press	press,
psykosen	psychosis,the psychosis,
georges	georges,
budet	the bid,the commandment,
miami	miami,
djupa	deep,
huruvida	whether,
sälja	sell,
finansieras	financed,funded,
djupt	deep,
säkra	reliable,safe,
serbiska	serbian,
tjeckoslovakien	czechoslovakia,
handeln	trade,
bibliska	biblican,biblical,
efterfrågan	demand,
gäst	guest,
export	export,
hittade	found,
skandinavien	scandinavia,
använts	was used,used,
genomsnitt	average,
planering	planning,
gammalt	old,
tvfilm	tv movie,
undviker	avoid,
klassificera	classifying,classify,
setts	observed,seen,
mankell	mankell,
stieg	stieg,
låten	the song,song,
sjunker	sinks,
markera	mark,
utsöndras	exudes,secreted,
uppvärmning	heating,warming,
mitt	my,center,
slut	end,out,
dateras	dated,
sommarspelen	summer games,summer olympics,
lång	long,
ljung	heather,
låna	borrow,
pressfrihetsindex	press freedom index,
substantiv	noun,
tillräcklig	sufficient,enough,
överlevde	survived,
bestämma	determining,decide,
oberoende	independent,
avsnittet	episode,
saken	the thing,matter,
saker	things,items,
förekommande	occuring,where,
mäta	compare,
främre	forward,front,
egna	own,
floder	rivers,
stanna	stop,
avrättade	executed,
tillbringade	spent,
mäts	is measured,
sektorn	sector,the sector,
floden	river,the river,
vidta	take,
stressorer	stressors,
glukos	glucose,
folkpartiet	liberal party,
konstruktion	construction,structure,
födelsetal	birthrate,birth rate,
val	choice,
idén	the idea,idea,
vad	as,
smeknamnet	nickname,
mäter	measuring,measure,
regisserad	directed,
vacker	beautiful,
nordamerikanska	north american,
lundell	lundell,
granne	neighbor,
hundratal	hundred,
ingått	entered,
stadens	the town's,the citys,
karta	map,
made	made,
rybak	rybak,
arne	arne,
tema	theme,
missnöjet	grievance,discontent,
jenny	jenny,
reaktorn	reactor,
problemet	the problem,
stormakter	world powers,great power,superpowers,
eu	eu,
utöva	exercise,
runor	runes,
kant	kant,
året	the year,years,
illinois	illinois,
book	book,
ursprunget	origin,
åren	the years,years,
intresse	interest,
juni	june,
behandlar	treat,
tolkas	is interpreted,interpretation,interpret,
tolkar	interprets,
shakespeares	shakespeare,
risker	risker,
personligen	individual,personally,
fira	celebrate,
ställningar	positions,
margaret	margaret,
markant	considerably,markedly,
risken	the risk,
cliff	cliff,
nödvändigtvis	by necessity,necessarily,
knappast	dead,
inledning	introduction,
bysantinska	byzantine,
simpson	simpson,
tidning	newspaper,
