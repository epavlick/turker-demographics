foster	embryo,fetus
schack	chess
loggbok	logbook,journal
stätta	stiles,tile,stile,ladder
resurs	resource
monografi	monografia,monography,monograph
koprolali	coprolalia
mullusfiskar	perch fish,goatfish
kvast	broom
sugga	soe,sow
mellanfot	metatarsus,metatarsal,metatarsal bones
fagocyt	phagocyte
draperi	curtian,curtain,drapery,daperi
reologi	rheology,reology
fotbeklädnad	footwear
ökenråttor	gerbil,gherbils,okenrattor,desert rats,gerbils
reduktion	reduction
rubrik	headline
peang	hemostat
azidgrupp	azide group,azide,azid group
ödleblad	lizard tail,houttuynia,chameleon plant
sats	clause,theorem; sets,statements,kit
befruktning	impregnation,fertilisation,insemination,fertilization
makadam	tarmac,crushed rock,macadam
flicka	girl
fåfotingar	pauropoda
spindlingar	cortinariaceae,cortinarius,fungal genus
väska	bag,leather case
fritid	free time,leisure time,freetime,leisure
bioetik	bioethic,bioethics
höftledsgrop	acetabulum,hip bone
neologi	neology,a new logical
långbåge	longbow,long bow,langbage
akondroplasi	achondroplasia,kondroplasia,akondroplasia
brushane	bird,ruff
antropogen	created by humans,an anthropogenic,antropog,antropogenic,anthropogenic
häcklöpning	hurdles,hurdling,hurdle race
stolpiller	suppository,suppositories,stolpills
gom	palate,mouth,roof of mouth
frekvens	frequencies,frequency
geomorfologi	geomorphology
ingenjör	engineering,engineer
producent	prodcuer,producer
depolarisering	depolarization
maffia	mob,mafia
fröväxter	spermatophyte,seed-bearing plants,seed plants,seed plant
laryngoskop	laryngoscopy,laryngoskop,laryngoscope
georgier	georgian,georgians
biogeografi	biogeography
likör	cordial,liqueur,liqeur,liquor,liquer
privilegium	privilege,prerogative
rede	nest,network
rorsman	helmsman,steersman
motorväg	freeway,motorway,highway,interstate
metionin	methione,methionine
högtryck	anticyclone
kupol	cupola,dome
kampanil	bell tower,bellfry; bell tower,campanile
giftsnokar	elapidae,poisonous snakes,elapids
zirkon	zirkon,zirconium,zircon
konsubstantiation	consubstantiation
hällristning	petroglyph,rock carvings,rock carving
ängssyra	sorrel
klimatologi	climatology,klimatologia
plattform	platform,platform, pad, rig
gräslök	chives
besserwisser	wiseacre,know-it-all,know-all,know it all,besserwisser
nätvingar	night wings,neuropterans,net-winged insects,neuroptera
baptism	baptist faith,baptist,baptism,baptists,bapist faith
havskattfiskar	goatfish,sea wolfs,catfish fishing,catfished,catfish,wolffish
bläckpenna	pen,quill
promemoria	memo,memorandum
