konsumtion	consumption,
okänd	unknown,
brevet	the letter,
nordisk	nordic,
reidar	reidar,
antisemitiska	antisemetic,
buddy	buddy,
likaså	also,
paris	paris,
spel	game,
edward	edward,
slå	hit,
albumen	the albums,
bli	become,
kommersiella	commercial,
passagerare	passenger,
mördade	murdered,
ägande	owning,
upptar	occupies,
stormaktstiden	great power period,
skicklig	skillful,
jack	jack,
försöka	try,
haber	haber,
chokladen	the chocolate,
venus	venus,
upp	up,
verklig	real,
rollfigurer	roll model,
horn	horns,
manus	script,
dennes	his,
ungerns	hungrarys,
avfall	waste,
upprätthåller	maintains,
tänkte	thought,
trodde	thought,
aktiva	active,
bidrar	contributes,
petra	petra,
med	with,
språken	languages,
prata	talk,
medelhavsklimat	mediterranean climate,
men	but,
hårda	hard,
drev	drove,
biografi	biography,
filosofen	the philosopher,
rysk	russian,
mer	more,
regnskog	rain forest,
herr	mister,
sidan	side,
bipolär	bipolar,
regerande	ruling,
geografiskt	geographically,
demokratier	democracies,
förblir	remains,
stoft	dust,
magnusson	magnusson,
isen	the ice,
systematiska	systematical,
biskop	bishop,
efterföljare	following,
strax	soon,
underliggande	underlying,
bro	bridge,
ansluta	connect,
total	total,
eftervärlden	the world,
bra	good,
stått	stood,
domare	judge,
skicka	send,
hörn	corner,
fotbollslandslag	national football team,
behandlingar	treatments,
supportrar	supporters,
återstående	remaining,
mercurys	mercurys,
övertala	convince,
holm	holm,
ansökte	applied,
wikipedias	wikipedias,
fermentering	fermentation,
köln	köln,
henri	henri,
kapitalistiska	capitalistic,
antiken	the ancient world,
mr	mr,
ofta	often,
sundsvall	sundsvall,
vietnamesiska	vietnamese,
partiets	parties,
vännen	the friend,
våldsam	violent,
utlöste	triggered,
befolkningsutveckling	population development,
vågen	the wave,
förväntade	expected,
talets	the speechs,
krävs	needs,
konstitutionen	constitution,
indier	indians,
polen	poland,
fröken	miss,
enhet	entity,
vänster	left,
nobelstiftelsen	nobel foundation,
kallare	colder,
trött	tired,
gillar	likes,
hos	with,
polis	police,
gata	street,
elektriskt	electric,
typen	the type,
biografer	movie theaters,
inrikes	domestic,
orsakar	causes,
åstadkomma	create,
neutralt	neutral,
förståelse	understanding,
barbro	barbro,
orsakat	caused,
sedd	seen,
klarar	do,
turkiet	turkey,
typer	types,
indelat	split,
orden	the words,
danny	danny,
medföra	result,
själva	self,
medlemsstat	member state,
grekiska	greek,
lämningar	remnants,
indelad	divided,
kända	known,
kontrollen	the control,
existera	exist,
arbetat	worked,
över	over,
arbetar	works,
kvicksilver	mercury,
förfäder	ancestors,
vart	each,
varv	dockyard,
ormar	snakes,
kampen	fight,
ibrahimović	ibrahimovic,
munnen	the mouth,
murray	murray,
varg	wolf,
besittningar	holdings,
buddhister	buddhists,
publicerade	published,
brinner	on fire,
nationell	national,
personal	staff,
friska	fresh,
infektioner	infections,
blott	merely,
upptagen	occupied,
band	band,
spelningen	the gig,
sverige	sweden,
hänga	hang,
avskaffandet	abolishment,
silver	silver,
jämförelser	comparison,
utvecklar	develops,
huvudartikel	main article,
debut	debut,
utveckling	development,
tillgängligt	available,
detroit	detroit,
diskuteras	discussed,
utvecklad	developed,
newport	newport,
angola	angola,
päls	fur,
germanska	germanian,
medier	media,
kontroverser	controversies,
serien	the series,
håret	the hair,
god	good,
hänvisa	refer,
ammoniak	ammonia,
ihop	together,
förändringar	changes,
behöva	need,
brukar	usually,
nationalistiska	nationalistic,
standard	standard,
neutroner	neutrons,
normer	standards,
anarkister	anarchists,
underordnade	subordinates,
statsministern	head of state,
väldiga	immense,
bredvid	next to,
vetenskapliga	scientific,
samhälle	society,
att	that,
befolkade	populated,
sökte	searched,
professionell	professional,
nyheter	news,
gå	go,
jamaica	jamaica,
sexuellt	sexual,
östberg	Östberg,
tecknade	drew,
leddes	was led,
sexuella	sexual,
tung	heavy,
begränsat	limited,
förklarade	explained,
xis	the eleventh's,
master	master,
punkter	points,
objekten	the objects,
hollywood	hollywood,
bitter	bitter,
tog	took,
adjektiv	adjective,
besegrades	defeated,
albert	albert,
kvarvarande	remaining,
skildes	was seperated,
meddelande	message,
roms	romes,
påverkad	influenced,
leden	the route,
formell	formal,
upphov	source,
sonen	the son,
slutsats	conclusion,
mjölk	milk,
trey	trey,
sheen	sheen,
utformningen	the layout,
tretton	thirteen,
obligatorisk	mandatory,
försörja	support,
nedgång	fall,
låta	let,
boston	boston,
filosofisk	philosophic,
rör	touches,
joakim	joakim,
växer	grows,
trakten	region,
omvandling	transformation,
industriellt	industrial,
lämnar	leaves,
lämnat	left,
situationer	situations,
magnus	magnus,
sjukvård	healthcare,
lades	put,
ulrich	ulrich,
anatomi	anatomy,
verkat	worked,
dessa	these,
flygplatser	airports,
bedrivs	conducted,
konserthus	concert hall,
utställning	exhibition,
fjädrar	feathers,
diskuterats	discussed,
övertog	overtook,
singer	singer,
arkitektur	architecture,
dom	conviction,
professor	professor,
dog	died,
metan	methane,
förlorar	loses,
grovt	heavy,
singel	single,
flod	river,
idrott	sports,
mitten	middle,
åsikten	the opinion,
hjälper	helps,
hus	house,
skyldig	responsible,guilty,
höjdpunkt	high point,
legitimitet	legitimacy,
senare	later,
rankning	ranking,
absolut	absolute,
sätter	puts,
tortyr	torture,
krönika	chronicle,
anländer	arrives,
buss	bus,
vinna	win,
ägare	owner,
rico	rico,
målvakt	goalee,
gods	domain,
lastbilar	truck,
kontinuerlig	continuous,
stycke	piece,
dj	dj,
tillståndet	the state,
de	the,
dygn	day,
kommunisterna	the communists,
samfund	order,
gogh	gogh,
stod	stood,
bensin	gasoline,
offret	the victim,
bas	base,
sköta	operate,
domaren	the judge,
konst	art,
utgåvan	the edition,
ursäkt	excuse,
tyngre	heavier,
fågelarter	species of bird,
lasse	lasse,
sutra	sutra,
publicerades	published,
blev	became,
tidningen	the newspaper,
kurdiska	kurdish,
zonen	the zone,
grundarna	founders,
historiens	historys,
gunnar	gunnar,
hamnar	lands,
öppnade	opened,
premiärminister	prime minister,
hedersdoktor	honorary degree,
allra	most,
materialet	material,
tanken	idea,
göta	göta,
rörelsens	movements,
israelisk	israeli,
intog	seized,
ber	asks,
maniska	manic,
kämpa	fight,
tilldelades	awarded,
världsturné	world tour,
schweiz	switzerland,
garanterar	ensures,
fns	un's,
tillämpas	applied,
beck	beck,
näringslivet	industrial life,
skalv	quake,
brad	brad,
anordnas	arranged,
nordiskt	nordic,
genus	genus,
graviditeten	the pregnancy,
verka	operate,
atombomberna	the nuclear bombs,
aktuell	current,
igelkotten	the hedgehog,
kännetecken	distinction,
tusentals	thousands,
räcker	enough,
uttalat	outspoken,
omstritt	controversial,
japans	japans,
fri	free,
socialistiskt	socialistic,
framträdande	apperance,
möjliggjorde	allowed,
frisk	healthy,
arbetslösheten	unemployment,
verktyg	tools,
barndom	childhood,
diktatorn	the dictator,
hitlers	hitlers,
tillämpa	administer,
omfatta	cover,
öster	east,
igång	start,
närvarande	present,
fest	party,
juridik	law,
spritt	spread,
kometer	comets,
chile	chile,
förstnämnda	first named,
vagn	carrige,
parterna	parties,
intag	intake,
slutliga	evenutal,
frankrikes	frances,
petrus	petrus,
tintin	tintin,
nationer	nations,
blåser	blowing,
sushi	sushi,
gärna	readily,
tänkare	thinker,
brittiskt	british,
sommar	summer,
madonna	madonna,
tät	compact,
påverkades	was affected by,
vänstern	western,
sagor	fairytales,
patent	patent,
bella	bella,
kommunistpartiets	the communist party,
utgivna	published,
äger	owns,
makt	power,
benämningar	terms,
djupare	deeper,
andelen	the share,
ökade	increased,
welsh	welsh,
funktionen	the function,
formatet	the format,
delstaten	the state,
yngsta	youngest,
bilen	the car,
återvända	return,
perspektiv	perspective,
finska	finnish,
nedan	below,
vetenskaplig	scientific,
charlie	charlie,
kampanj	campaign,
dåvarande	formerly,
mamma	mother,
roma	roma,
jean	jean,
fortplantning	reproduction,
kraftigt	heavily,
gärningsmannen	culprit,
newton	newton,
dödsoffer	casualty,death victim,
norsk	norwegian,
körs	being driven,
bollen	the ball,
grader	degrees,
utrotning	extinction,
beskriver	describes,
kroppens	the bodies,
döda	dead,
kalender	calender,
kolväten	the hydrocarbon,
matteus	matteus,
använt	used,
distributioner	distributions,
huvud	head,
lunginflammation	pneumonia,
borgen	the castle,
hav	seas,ocean,
maya	maya,
återgick	returned,returning,
everton	everton,
engelskans	english,
uppmärksammade	observed,
hepatit	heptatitis,
årlig	yearly,
modersmål	native language,
konsert	concert,
gandhi	gandhi,
hund	dog,
gifter	marries,
litauen	lithuania,
transkription	transcript,
kemiska	chemical,
sixx	sixx,
kunna	be able,
befolkningen	the population,
släkt	family,
befann	located,
borg	tower,castle,
delade	split,
humor	humour,
varierande	varying,
beroendeframkallande	addictive,
miljöproblem	environmental problems,
princip	principle,
akademi	academy,
säsongerna	seasons,
shakespeare	shakespeare,
utse	name,
litterära	literal,
karaktäriseras	characterizes,
deltagarna	participants,
annan	another,
stadsdelarna	districts,
monoteism	monotheism,
ishockeyspelare	ice hockey player,
burj	burj,
hörde	heard,
vägar	roads,
olympiska	olympic,
bolt	bolt,
möjligheterna	the possibilities,
hotellet	the hotel,
meyer	meyer,
fördelen	the advantage,
förslaget	the suggestion,
mycket	much,
tillverkas	manufacture,
strömmar	streams,
förknippade	associated,
olika	different,
förgäves	in vain,
jacques	jacques,
tydliga	obvious,
hänt	happened,
återfinns	is rediscovered,
grundades	was founded,
delvis	partially,
marshall	marshall,
som	which,
menade	meant,
tydligt	obvious,
spåra	track,
varmare	warmer,
lagt	laid,
kjell	kjell,
nova	nova,
fria	free,
gia	gia,
förebild	role model,
etablerat	established,
fadern	the father,
skulden	the guilt,
själv	alone,
offer	victim,
trenden	the trend,
berg	mountain,
verde	verde,
tigern	the tiger,
skulder	debts,
avsevärt	substantially,
definierade	defined,
partiledare	party leader,
drabbat	affected,
gymnasiet	high school,
emil	emil,
polska	polish,
studierna	the studies,
slaviska	slavic,
litterär	literary,
långvarig	long,
pest	plague,
regeringen	the government,
driva	operate,
tillika	also,
araber	arabs,
avsnitt	episode,
föregångare	predecessor,
xiis	xii,
handelspartner	trading partner,
krävde	demanded,
empati	empathy,
publiceringen	publishing,
liberalism	liberalism,
handel	trade,
förmåga	ability,
möte	meeting,
dotter	daughter,
tim	tim,
arkitekter	architects,
digital	digital,
möts	meets,
nr	number,
götaland	götaland,
mexikanska	mexican,
avskaffades	was abolished,
femton	fifteen,
bostadsområden	residential areas,
vintrarna	the winters,
modell	model,
tävling	competition,
jehovas	jehovas,
reglerar	regulates,
rött	red,
totalt	complete,
vagnar	carriges,
trettio	thirty,
långtgående	far-reaching,
bergmans	bergmans,
funktionerna	the functions,
bomben	the bomb,
uppfanns	invented,
global	global,
datum	date,
uppgifter	tasks,
tredje	third,
stödjer	supports,
bomber	bombs,
inkomst	income,
machu	machu,
vikingarna	the vikings,
religion	religion,
mottagarens	the reciever,
fängelset	prison,
dä	the elder,
då	then,
intresserade	interested,
petersburg	petersburg,
vem	who,
musikstilar	music genres,
serbiens	serbias,
fördrevs	was banished,
lättare	easier,
varvid	in which,
kompositörer	compositors,
krossa	crush,
metod	method,
sätt	way,
afrikansk	african,
olyckor	accidents,
levnadsstandard	standard of living,
olympia	olympia,
idéer	ideas,
heinz	heinz,
jämnt	evenly,
villa	house,
trend	trend,
reklamen	the commercial,
stilar	styles,
jämna	even,
rymden	space,
svartån	svartån,
utlösning	ejaculation,
hästen	the horse,
bakom	behind,
firandet	the celebration,
stimulera	stimulate,
måne	moon,
södra	south,
kunskapen	the knowledge,
utspelar	takes place,set,
somalia	somalia,
kön	gender,
gräs	grass,
gazaremsan	the gaza strip,
köket	the kitchen,
kärlek	love,
påstår	claims,
oerhört	tremendously,
katten	the cat,
beskrivits	described,
versioner	versions,
antarktiska	antarctic,
bor	lives,
kemi	chemistry,
bärande	leading,
mellankrigstiden	interwar years,
franklin	franklin,
tilltagande	increasing,
mänsklighetens	humanities,
studier	studies,
diagnosen	diagnosis,
dåtidens	past times,that time,
burr	burr,
vapnet	the weapon,
utövas	is practised,
världshälsoorganisationen	world health organization,
basen	became,
biträdande	assisting,
förteckning	listing,
modellen	the model,
trinidad	trinidad,
kärnkraftverk	nuclear power plant,
sprids	spreads,
abstrakta	abstract,
ande	spirit,
inblandade	involved,
emellan	between,
regel	rule,
kristian	kristian,
grundläggande	primary,
förbjöds	forbidden,
ställt	taken,put,
fransmännen	the french,
typerna	the types,
relationerna	the relationships,
övergå	transend,
målvakten	the goalkeeper,
närmar	closing,
norrköpings	norrköpings,
styras	steered,
fly	escape,
löner	salaries,
ibm	ibm,
tokyo	tokyo,
läkemedel	medicine,
partnern	the partner,
mästarna	the champions,
interaktion	interaction,
frukt	fruit,
kombination	combination,
vittnen	witnesses,
domkyrka	cathedral,abbey,
bristande	wanting,lack,
generell	general,
erbjuder	offers,
ulf	ulf,
hiroshima	hiroshima,
några	a few,
december	december,
winston	winston,
gentemot	towards,against,
abort	abortion,
hemliga	secret,
dennis	dennis,
genomgått	experienced,
milda	mild,
oslo	oslo,
engelsmännen	the british,
ekonomiska	economical,
begick	commited,
simning	swimming,
muslimerna	the muslims,
nikolaj	nikolaj,
industriell	industrial,
perserna	the persians,
regeringstid	term of government,
överensstämmer	conform,
fascism	fascism,
utlandet	abroad,
familjens	the familys,
nyligen	recently,
läkare	doctor,
göteborgs	gothenburgs,
maj	may,
mao	mao,
asien	asia,
bergarter	rock types,
stöds	is supported,
flyttas	moved,
benny	benny,
tala	speak,
basket	basketball,
sa	said,
ida	ida,
vintrar	winters,
komplicerad	complicated,
landshövding	county governor,
ganska	quite,
unionen	the union,
huvudsak	main thing,
generalguvernören	general governor,
motståndet	the resistence,
böcker	books,
verksam	active,
landskap	province,
linköping	linköping,
organisation	organization,
jim	jim,
tilldelats	awarded,
behandlingen	the treatment,the treament,
sekter	sects,
äkta	genuine,
nazisterna	nazis,
försvaret	the defense,
växte	grew,
öppnades	was opened,
halt	stop,
janeiro	janeiro,
domstolar	courts,
matcher	games,
författarna	writers,
komponenter	components,
hamilton	hamilton,
matchen	the game,
kantoner	cantons,
färgen	the color,
vindkraft	wind power,
organ	body,
växa	grow,
opera	opera,
förväxlas	confused,
omöjligt	impossible,
stockholm	stockholm,
hotad	threatened,
dominerar	dominates,
runstenar	runestones,
bildning	education,form,
tysklands	germanys,
födelsedag	birthday,
en	a,
stående	standing,
citat	quote,
ed	ed,
utbrett	wide,
står	standing,
vattendrag	streams,
avkomma	offspring,
resultera	result,
ledamöter	commissioners,
kött	meat,
er	you,
album	album,
teorier	theories,
medelhavsområdet	the mediterranean area,
bly	led,
stortorget	stortorget,
sjuka	sick,
accepterar	accepts,
pamela	pamela,
områdena	the areas,
tronföljare	successor,
kattdjur	cat,
metro	metro,
våra	our,
bytt	traded,
juldagen	christmas day,
zuckerberg	zuckerberg,
välkänd	well known,
byta	trade,
pund	pound,
politiker	politician,
självmord	suicide,
traditioner	traditions,
rankningar	rankings,
gordon	gordon,
processen	the process,
kommentar	comment,
laboratorium	laboratory,
origin	origin,
xi	xi,
här	here,
hård	hard,
begår	commits,
akademien	academy,
centralt	central,
skapandet	the making,
hårt	hard,
okända	unknown,
teologi	teology,theology,
består	exists,
grundämnen	elements,
desmond	desmond,
nästa	next,
williams	williams,
vilka	who,
anus	ass,
kronprinsessan	crown princess,
färre	less,
kallade	called,
fysiskt	physical,
irakiska	iraqi,
tillräckliga	insufficient,sufficient,
svenskarna	the swedes,
bönder	farmers,
provins	province,
beslutet	the decision,
smeknamn	nickname,
europeisk	european,
passade	suiting,
marinen	navy,
genomsnittet	average,
framställning	production,
sidorna	the pages,pages,
kamprad	kamprad,
motståndarna	the opponents,
medlemmarna	the members,
ändrades	changed,
modeller	models,
fordon	vehicle,
afrikanska	african,
tiotusentals	tens of thousands,
kromosomerna	the chromosomes,
konsekvenser	consequences,
församlingar	parishs,
grundar	bases,
jordskorpan	earth crust,
allen	allen,
västberlin	west berlin,
kevin	kevin,
medvetande	consciousness,
priserna	the prices,
hjälp	help,
nikola	nikola,
explosionen	the explosion,
förste	the first,
zon	zone,
etiopiska	ethiopian,
centralbanken	central bank,
förhållandena	conditions,
gustavs	gustavs,
kust	coast,
finlands	finlands,
norman	norman,
knutna	associated,
religionen	the religion,
betyda	mean,
politisk	political,
dvärgar	dwarfs,
glödlampor	light bulbs,
america	america,
 miljoner	millions,
civilisationer	civilizations,
lyfter	lifts,
norrmän	norwegians,
varken	either,
täcks	covers,
öppet	open,
ursprung	root,
fredspriset	peace prize,
nordligaste	northern,
runda	round,
drivs	driven,
engagemang	commitment,
herren	the lord,
marocko	marocco,
japansk	japanese,
perfekt	perfect,
tror	believe,
bandets	the bands,
rötter	roots,
guld	gold,
motivet	the motive,
passande	fitting,suitable,matching,
historien	history,
statsmakten	power,
hockey	ice hockey,
sierra	sierra,
ovanliga	unusual,
ges	be given,
jazz	jazz,
folkomröstning	referendum,
platta	flat,
facupen	fa-cup,
undersöka	research,
rasen	the race,
drabbar	troubles,
påminner	reminds,
reser	travels,
ländernas	the countries,
artist	artist,
skivkontrakt	record contract,
råd	council,
dianno	dianno,
spridda	spread,
vara	be,
erbjöds	offered,
minnen	memories,
underlätta	ease,
brännvin	schnaps,
snabbare	faster,
terräng	terrain,
teoretisk	theoretical,
skärgård	archipelago,
talman	spokesperson,
stanley	stanley,
sport	sport,
menar	means,
kandidater	candidates,
enhetlig	uniform,
försvarsmakten	national defense,
katastrofer	catastrophes,
kritiserade	critisized,
begränsningar	limitations,
konstaterade	established,
kilometer	kilometer,kilometers,
önskade	wished,
import	import,
kommunismens	the communisms,
katastrofen	the catastrophy,
yta	surface,
återigen	yet again,
anledningarna	the reasons,
hämtat	collected,
utgivningen	the publication,
konstnären	the artist,
jr	junior,
åker	go,
glenn	glenn,
timme	hour,
bekämpa	fight,
amerikanska	american,
dödade	killed,
uppskattade	appreciated,
kirsten	kirsten,
warhol	warhol,
spelfilmer	motion pictures,
ordagrant	literal,
engagerade	engaged,
spindlar	spiders,
ståndpunkt	standpoint,
år	year,
nils	nils,
benämningen	the name,
gjorde	did,
placerar	places,
tum	inch,
pakistan	pakistan,
vilja	will,
statschefen	the head of state,
pop	pop,
termen	the term,
statsreligion	state religion,
hamnade	landed,
östtyska	east german,
uppehåll	hiatus,
handlande	action,
drogs	was pulled,
skånska	scanian,
mätningar	measurements,measurments,
långfilm	feature film,
lexikon	lexicon,
barry	barry,
förekomsten	presence,
mark	ground,
oden	oden,
lidit	suffered,
hämtade	brought,
knappt	barely,
socialdemokrater	social democrats,
mary	mary,
kultur	culture,
dräkt	costume,
anderna	the andes,
partido	partido,
bmi	bmi,
använder	uses,
bilderna	the pictures,
prinsessan	the princess,
fiende	enemy,
uppstod	developed,
situation	situation,
ansikte	face,
pippi	pippi,
insåg	realized,
kenya	kenya,
blad	leaves,
beteckna	denote,
grönland	greenland,
programvara	software,
världsbanken	world bank,
paz	paz,
försäkra	make sure,
långa	long,
ärftliga	genetic,
träffar	meets,
samt	also,as well as,
singapore	singapore,
skivbolaget	record label,
älskar	loves,
protoner	protons,
persons	persons,
målningar	paintings,
linjerna	the lines,
privilegier	privileges,
producerad	produced,
tradition	tradition,
fredspris	peace prize,
aktuella	current,
moder	mother,
kommunistisk	communistic,communist,
breda	wide,
avses	regard,
mynning	outfall,mouth,
medellivslängd	average lifespan,
nicklas	nicklas,
skandinaviska	scandinavic,
summer	sommar,
kommentarer	comments,
koncentration	concentration,
familjer	families,
harrison	harrison,
moçambique	mozambique,
reaktioner	reactions,
resa	travel,
libyen	libya,
ideologiskt	ideological,
utvinns	extracted,
rose	rose,
transeuropeiska	transeuropean,
lagerkvist	lagerkvist,
rosa	pink,
miljon	million,
gotland	gotland,
ideologiska	ideological,
nazismen	nazism,
infördes	introduced,
euron	the euro,
trä	wood,
guldbollen	guldbollen,
slöts	signed,
irland	ireland,
marcus	marcus,
sköttes	operated,
stund	while,
östergötland	Östergötland,
utrikespolitik	foreign affairs,
prägel	mark,
tillbehör	accessory,
amy	amy,
test	test,
vampyrer	vampires,
klimat	climate,
mod	courage,
afrikas	africas,
skadade	wounded,
adams	adams,
republik	republic,
födde	gave birth too,
gröna	green,
intet	nothing,
nämnas	mentioned,
skyddar	protects,
innebära	mean,
monopol	monopoly,
huvudrollen	leading part,
eddie	eddie,
gång	time,
lågt	low,
präglades	imprinted,
alkoholer	alcohols,
verksamheter	operations,
strindberg	strindberg,
maos	mao's,
jordbruket	the agriculture,
slår	beats,
slås	is hit,
fört	lead,
konsten	the art,
buddha	buddha,
berodde	depended,
tunnlar	tunnels,
londons	london's,
olof	olof,
utskott	organ,
geografi	geography,
jacksons	jacksons,
oliver	olives,
kaffet	the coffee,
tyske	german,
ideologi	ideology,
om	if,
indianska	native american,
herrlandslag	men's national team,
sri	sri,
populationen	the population,population,
metaforer	metaphores,
lyssnade	listened,
förbundskapten	manager,
bidragen	contributions,
spelen	the games,
visst	certain,
befäl	command,
berger	berger,
lands	on land,
lagarna	the laws,
partiet	the party,
klassiker	classic,
nådde	reached,
överföras	transferred,
karriär	career,
intellektuella	intellectuals,
gravid	pregnant,
behandling	treatment,
stark	strong,
evangeliska	evangelical,
start	start,
anställd	hired,
specifika	specific,
talades	spoke,
gånger	times,
närmaste	closest,
fastställa	confirm,
rockband	rock band,
mars	march,
jul	christmas,
inriktning	direction,orientation,
land	country,
sämsta	worst,
bevarad	kept,
gången	time,
egen	own,
traditionerna	the traditions,
minne	memory,
ekonomi	economy,
jamaicas	jamaicas,
kvartsfinalen	quarter finals,
minns	remembers,
vinkeln	the angle,
kröntes	crowned,
kostar	costs,
ac	ac,
följde	followed,
gustafs	gustafs,
youtube	youtube,
närmast	closest,
fjorton	fourteen,
öns	the islands,
bronsåldern	the bronze age,
pontus	pontus,
godkände	approved,
knut	knot,
asteroider	astroids,
blues	blues,
vanliga	regular,usual,
ökande	increasing,
rubiks	rubik's,
många	many,
omgivande	surrounding,surounding,
stannade	stayed,
avslöjade	revealed,
genren	genre,
däremot	on the contrary,
koppar	copper,
gifte	married,
kvarstod	remained,
rykten	rumors,
erövring	conquest,
missbruk	abuse,
medverkar	contributes,contribute,
världsliga	worldly,
kväll	evening,
skuggan	the shadow,
morgonen	the morning,
vinner	wins,
beteckning	label,
därvid	therewith,
snabbaste	fastest,
decennierna	decades,
resolution	resolution,
renässans	renaissance,
olympiastadion	olympa stadium,
vila	rest,
släppt	released,
alf	alf,
separat	seperate,
öknen	the desert,desert,
konsekvent	consistent,
kammare	chamber,
samhällen	communities,
spelade	played,
levern	the liver,
atlanta	atlanta,
zink	zinc,
skogarna	the forests,
påbörjades	was started,
röstade	voted,
symboler	symbols,
kasta	throw,
ansluter	connects,
fas	phase,
avhandling	thesis,
får	can,
israeliska	isrealic,
strand	beach,
kulminerade	culminated,
unionens	the union's,
tjeckiska	czech,
djurarter	species,
knutsson	knutsson,
louis	louis,
muslimska	muslim,
harry	harry,
rod	rod,
medel	middle,
döttrar	daughters,
grekland	greece,
påståenden	claims,
egendom	property,
dödsstraff	death penalty,
utökade	expanded,
utåt	outwardly,
givaren	the giver,
tvskådespelare	tv actor,
bedrev	managed,
stängt	closed,
publik	audience,
misstänkta	suspected,
islams	islams,islam's,
hänsyn	consideration,
gruppen	the group,
upptäcka	discover,
kronor	kronor,
observeras	observed,
grupper	groups,
lämna	leave,
jackie	jackie,
boxning	boxing,
exklusiv	exclusive,
kärnvapen	nuclear weapons,
våg	road,
traditionellt	traditional,
hoppades	hoped,
social	social,
oftare	more often,
tillkännagav	announced,
varelser	creatures,
medlemskap	membership,
samlade	collected,
nazityskland	nazi germany,
ordinarie	regular,
vin	wine,
grunda	found,
kritiserat	criticised,
dahlén	dahlén,
enat	united,
främja	further,
biskopen	the bishop,
sitter	sit,
representeras	represented,
representerar	represents,
dödligt	deadly,
torra	dry,
reptiler	reptiles,
permanenta	permanent,
cellerna	the cells,
akademiens	the academy's,
berättade	told,
romersk	roman,
vm	world championship,
koma	coma,
räknar	counts,
graven	the grave,grave,
lagstiftande	legislating,
bror	brother,
undergång	doom,
östra	eastern,
investeringar	investments,
flytt	escaped,
tillverkningen	production,the production,
kryddor	spices,
sociala	social,
kapitalism	capitalism,
läkaren	the doctor,
jakob	jakob,
nordvästra	north western,
bosatt	resident,
betoning	stress,
medförde	resulted,brought,
födseln	the birth,
järnvägsnätet	railroad network,
historiskt	historic,historical,
vägnätet	road network,
hugo	hugo,
faktum	fact,
försvinner	disappears,
uttrycka	express,
reidars	reidars,
makter	powers,
hoppade	jumped,
variant	variety,
betraktades	regarded,
pettersson	pettersson,
grundämne	element,
fötts	born,
vattenkraft	hydroelectric power,
praktiska	practical,
enzymer	enzymes,
anklagade	accused,
tsar	tsar,
homosexuella	homosexual,
rockgrupper	rock bands,
juan	juan,
civila	civil,
hållit	held,
september	september,
längd	length,
scott	scott,
vietnamkriget	vietnam war,
människans	humans,mankinds,
hundratusentals	hundreds of thousands,
humör	mood,
rike	kingdom,
alla	all,
rika	rich,
caesars	caesars,
miljön	the environment,
längden	lenght,
abbey	abbey,
systems	systems,
stadshus	town hall,
österrikes	austrias,
argentina	argentina,
gustafsson	gustafsson,
suverän	terrific,
offensiven	offensive,
beräkna	calculate,
elden	the fire,
petter	petter,
grekisk	greek,
producerat	produced,
introducerade	introduced,
producerade	produced,
olycka	accident,
försöken	the tries,
journalisten	the journalist,
fulla	complete,
namibia	namibia,
skrivit	written,
journalister	journalists,
genom	through,
kontinentens	the continents,
försöker	tries,trying,
ifk	ifk,
etnisk	ethnic,
enstaka	occasional,
england	england,
mental	mental,
positionen	the position,
betyg	grades,
fisk	fish,
flytta	move,
energi	energy,
mongoliet	mongolia,
ollonet	the glans,
oftast	most often,
kopplad	connected,
garvey	garvey,
infrastrukturen	infrastructure,
ölet	the beer,
forskning	research,
förföljelser	pursuits,persecutions,
rowling	rowling,
ingående	enter into,
lungorna	the lungs,
sparken	gets fired,
alltmer	more and more,
stöder	supporting,
stjärnor	stars,
ersatt	replaced,
knäppupp	knäppupp,
omfattande	large,
kostade	cost,
ökat	increased,
vasas	vasas,
trummisen	the drummer,
svarade	answered,
turistmål	tourist attraction,
stavningen	the spelling,
finland	finland,
skilja	seperate,
konsumtionen	consumption,
förkortning	abbreviation,
underhåll	allowance,
ytterligare	additional,
ensam	alone,
nivåer	levels,
besök	visit,
sändes	was sent,
etiska	ehtical,
bidragit	contributed,
arsenal	arsenal,
treenighetsläran	school of trinity,
minoritetsspråk	minority language,
spekulationer	speculations,
bland	including,
synes	appears,
rygg	back,
förbi	past,
kom	came,
liknas	compared to,
misslyckas	fails,
stort	big,
definitioner	definitions,
lördagen	the saturday,
storm	storm,
sår	wound,
växthusgaser	greenhouse gas,
luminositet	luminosity,
besläktat	related,
serotonin	serotonin,
triangeln	the triangle,
borgmästare	mayor,
två	two,
växterna	plants,
humanistiska	humanistic,
fred	peace,
obama	obama,
följden	result,
långsamt	slowly,
återkom	returned,
direkt	direct,
einsteins	einsteins,
andersson	andersson,
personens	the persons,
stjärnan	the star,
avtar	declines,
försökte	tried,
kusin	cousin,
avslutade	ended,
inkluderar	includes,
generationen	the generation,
tvärtom	on the contrary,
motsatte	opposed,
mountain	mountain,
visats	shown,
vägen	the road,
infrastruktur	infrastructure,
lik	alike,
caesar	caesar,
förmögenhet	wealth,
unga	young,
unge	kid,
världsarvslista	world heritage list,
krafter	forces,
gillade	liked,
stjärnans	the stars,
freddie	freddie,
sydostasien	south east asia,
dagligt	daily,
plan	level,
utbrott	outbreak,
utgör	constitutes,
organiserade	organized,
kombinationer	combinations,
sånger	songs,
arter	species,
forskarna	the scientists,
utsattes	subjected,
ko	cow,
km	kilometers,
kanalen	the channel,channel,
influensan	the influenza,
sången	the song,
organisk	organic,
mesopotamien	mesopotamia,
gudarna	the gods,
ingenting	nothing,
presidentens	the presidents,
detalj	detail,
kolonialism	colonialism,
antagit	presumed,
därifrån	from there,
undre	lower,
wallenberg	wallenberg,
beräkningar	calculations,
medverka	participate,
åländska	Åland swedish,
axel	axel,
jämfört	compared,
kontor	office,
inklusive	including,
vardera	each,
tekniker	technician,
typiska	typical,
husen	the houses,
skickas	is sent,
skickar	sends,
avsaknaden	absence,
tvkanaler	tv channels,
mediciner	medicines,
byter	exchanges,
tidszon	timezone,
norrköping	norrköping,
någon	someone,
kriterier	criteria,
etiopien	ethiopia,
maurice	maurice,
suveränitet	sovereignty,
vind	wind,
sex	six,
arg	angry,
järnväg	railway,
händelsen	the occurence,
mörkare	darker,
pär	pär,
guinea	guinea,
uppskatta	appreciate,
fission	fission,
jakten	the hunt,
alqaida	al-qaida,al-qaeda,
hellström	hellström,
champagne	champagne,
bildandet	establishment,
giftermål	marrige,
kategorin	the category,
rörelserna	the movements,
likhet	resemblance,
kritiserades	critisized,
revolutionen	the revolution,
stadsdel	district,
demografiska	demographical,
forskare	scientists,
bästa	best,
musklerna	the muscles,
tiderna	the times,
uppfattning	understanding,
stå	stand,
kamp	fight,
kyrkliga	religious,
globala	global,
hypotesen	the hypothesis,
kroatiens	croatias,
läsaren	the reader,
bell	bell,
betydde	meant,
sweet	söt,
tennessee	tennessee,
belägna	located,
hypoteser	hypothesis,
merparten	most,
kungafamiljen	the royal family,
johannes	johannes,
idén	the idea,idea,
oändligt	infinitely,
byxor	pants,
ska	will,
skönhet	beauty,
inför	before,
walter	walter,
östafrika	east africa,
bengt	bengt,
popularitet	popularity,
budgeten	the budget,
gas	gas,
togs	taken,
rak	straight,
anthony	anthony,
rättigheterna	the rights,
vann	won,
trupperna	troops,the troops,
detsamma	the same,
delades	split,
motorväg	highway,
framträder	appear,
socialism	socialism,
döptes	baptised,
hegel	hegel,
läser	read,
bestående	comprising,lasting,
radio	radio,
casino	casino,
inspelningar	recordings,
von	von,
ris	rice,
alaska	alaska,
legender	legends,
lokaler	place,
korruptionsindex	corruption index,
lagar	laws,
tillfällen	oppertunities,
kombineras	combined,
rederiet	shipping company,
staffan	staffan,
skeppen	the ships,
kombinerat	combined,
demografi	demographics,
möjlighet	oppertunity,
tidpunkten	the time,the moment,
listor	lists,
barnen	children,
kombinerad	combined,
administrationen	administration,
tyder	indicates,
spears	spears,
inledde	started,
laddning	charge,
sapiens	sapiens,
utmed	along,
kungahuset	royal house,
snarare	rather,
republiken	the republic,
berömt	praised,
debatten	the debate,
avlägsna	remove,
mot	against,
älska	love,
normala	normal,
albanien	albania,
jorderosion	earth erosion,
ministerrådet	minister counsellor,
normalt	normally,
person	person,
dikter	poems,
nutid	present,
präglad	marked,
följande	following,
kontakter	contact,
nacka	nacka,
stränder	beaches,
komplett	complete,
fredliga	peaceful,
remmer	remmer,
finansiella	financial,
tropisk	tropical,
fascistiska	fascistic,
festivalen	the festival,
administrativt	administrative,
skall	shall,
minoriteten	minority,
nordväst	north west,
festivaler	festivals,
åtal	prosecution,
strävan	the quest,
varuhus	department store,
djup	deep,
bestå	consists,exist,
producerats	produced,
synnerhet	specially,
gör	makes,
herre	lord,
enklare	simpler,
möttes	met,
bit	piece,
begravdes	buried,
användas	used,
kolonialtiden	the colonial times,
miami	miami,
arthur	arthur,
hittas	found,
minskning	decline,
begärde	demanded,
lindgrens	lindgrens,
möjlig	possible,
tolkats	interpreted,
byggnader	buildings,
egyptiska	egyptian,
saknas	missing,
våldet	the violence,
körberg	körberg,
krigare	warrior,
byggnaden	building,
cocacola	coca cola,
västergötland	västergötland,
sammanhängande	connective,
vilda	wild,
trafiken	the traffic,
bildar	form,
pratar	talks,talking,
anne	anne,
saab	saab,
säger	says,
höjder	heights,
lösningen	the solution,
därför	because,
steg	rose,
italienska	italian,
producent	producer,
sten	stone,
plocka	pick,
lånat	borrowed,
engelske	english,
judendom	judaism,
kinesisk	chinese,
bosättningar	settlements,
personen	the person,
övergick	transended,
gemenskaperna	community,
efterträdare	successor,
linjer	lines,
edvard	edvard,
länderna	the countries,
socialistisk	socialistic,
industrialiserade	industrialized,
inte	not,
lager	layer,
efterföljande	subsequent,
spridas	spread,
öl	beer,
snarast	as soon as possible,
popsångare	pop singer,
medborgarna	the citizens,
rammstein	rammstein,
semifinalen	semi finals,
seger	victory,
institut	institution,
sprida	spread,
fast	even though,
jugoslavien	yugoslavia,
visas	shown,
knuten	tied to,
jonsson	jonsson,
regionen	the region,
ledamot	representative,
fralagen	the fra law,
serie	cartoon,
atom	atom,
kritisk	critical,
regioner	regions,
junior	junior,
lina	lina,
fader	father,
turné	tour,
ute	out,
planeternas	the planets,planets,the planets',
ledningen	the lead,
högt	high,
ur	out,
smycken	jewlery,
malin	malin,
erövrades	concoured,
planer	plans,
guyana	guyana (name),
tolka	interpret,
passera	pass,
chelsea	chelsea,
öland	öland,
tidens	time's,
titel	title,
nämner	mentions,
förbjudna	forbidden,
avsåg	meant,
detaljer	details,
intressanta	interesting,
avsattes	dismissed,
hårdrock	hard rock,
igenom	through,
personlighetsstörning	personality disorder,
räkna	count,
voltaire	voltaire,
psykoterapi	psychotherapy,
nordafrika	north africa,
möter	meets,
matematiker	mathematician,
manhattan	manhattan,
berättar	tells,
förr	sooner,
korn	korn,
beräknar	values,
medina	medina,
drag	move,
ägnar	spend time,
matematiska	mathematical,
riskerar	risks,
användbara	usable,
tillfälligt	temporarly,temporary,
alltså	therefore,
oväntat	unexpected,
passagerarna	passengers,the passengers,
uppträdande	performance,conduct,
produkt	product,
tunga	tongue,
ställe	place,
judisk	jewish,
hertig	duke,
nasa	nasa,
nash	nash,
inspelning	recording,
persbrandt	persbrandt,
alltför	all too,
ställa	set,
ge	give,
go	go,
träd	tree,
kolonialismen	the colonialism,
världsrekord	world record,
intensivt	intensive,
simon	simon,
turkisk	turkish,
fortfarande	still,
sena	late,
tillhör	belongs,
protokoll	protocol,
varierar	varies,
georgien	georgia,
hustru	wife,
medverkade	participated,
epost	email,
kommunistiska	communistic,
avslutas	ends,
avslutat	completed,
historikern	historian,
kommunismen	communism,
tävlingar	competitions,
eva	eva,
joel	joel,
noter	notes,
utbredning	distrubution,
romerska	roman,
utanför	outside,
överlevt	survived,
min	my,
månens	the moons,
warszawa	warsaw,
joey	joey,
riktigt	real,
derivator	derivative,
åtta	eight,
honan	the female,
geologiska	geological,
influerad	influenced,
anderssons	anderssons,
motsättningar	oppositions,
påsken	easter,
mussolini	mossolini,
folk	people,
kinas	chinas,
sträcker	stretches,
går	goes,
assisterande	assisted,
chicago	chicago,
skrivna	written,
byttes	was exchanged,
indiens	indias,
suveräna	terrific,
gamle	old,
koloni	colony,
eminem	eminem,
åtgärder	measures,
definitionen	the definition,
astrid	astrid,
teater	theater,
honom	him,
svårigheter	difficulties,
ukraina	ukraine,
motorvägarna	the highways,
innehar	holds,
ep	ep,
elektronik	electronics,
titanic	titanic,
springsteens	springsteens,
katolicismen	catholisism,
lagförslag	bill,
opinion	opinion,
översättningar	translations,
privata	private,
stundom	somtimes,
zlatan	zlatan,
förlora	lose,
avsedda	intended,
nåd	mercy,grace,
anatolien	anatolia,
övergår	surpasses,
keramik	ceramics,
tar	takes,
usa	usa,
fel	errors,
fem	five,
hemlig	secret,
kunde	could,
söder	south,
oktober	october,
orkester	orchestra,
inlandet	inland,
konservatism	conservatism,
utropade	cried out,
samspel	teamwork,
självständighet	independence,
penis	penis,
invigningen	the opening,
huxley	huxley,
organisationen	the organization,
vägrade	refused,
tillräcklig	sufficient,enough,
reguljära	regular,
baserad	based,
automatiskt	automatic,
baseras	based on,
väldet	the rule,
titlar	titles,
ingå	be included in,
process	process,
liknade	looked like,
ledamöterna	commisioners,
mozarts	mozart's,
talat	spoke,
fett	fat,
sydöstra	south east,
talar	speaks,
saknade	missed,
lanserade	introduced,
övergrepp	assault,
brian	brian,
internationella	international,
undantaget	except,
folkmängd	population,
sin	its,
kriminella	criminal,
fara	danger,
väpnad	armed,
monica	monica,
billiga	cheap,
mötte	met,
spannmål	grain,
tack	thanks,
religiös	religious,
utfördes	preformed,
regeringsmakten	government power,
säljer	sells,
lundgren	lundgren,
drabbats	afflicted,
kommunikationer	communications,
kvinnliga	female,
handboll	handball,
fungerade	working,
presidenter	presidents,
plats	place,
universiteten	the universities,
hunnit	had time to,
cambridge	cambridge,
karlstad	karlstad,
blandas	mixes,
offentligt	publicly,
verklighet	reality,
listan	the list,
uppdelat	split,
egna	own,
tecknet	the sign,
tvungna	forced to,
uppdelad	split,
lärjungar	disciple,
insekter	insects,
referenser	references,
utfärdade	issued,
zagreb	capital of croatia,
fler	more,
ägna	spend,
periodiska	periodic,
intäkterna	the revenues,
runt	around,
sönder	broken,
delar	parts,
kläder	clothes,
beslut	decision,
förmågor	abilities,
växande	growing,
säsonger	seasons,
skog	wood,
humanism	humanism,
fortsätta	continue,
smallwood	smallwood,
populärmusik	popular music,
 procent	percent,
intresset	the interest,
säsongen	season,
banan	banana,
programmet	the application,
uppfattar	percieves,
endast	merely,
nödvändiga	essential,
kritik	critisism,
uggla	owl,
minskad	decreased,
hantverkare	handy worker,
samarbetat	collaborated,
kapitalismens	capitalism's,
max	max,
solsystem	solar system,
minskat	decreased,
plural	plural,
förutsättningar	condition,
hörs	heard,
egenskaperna	the qualities,
påverkats	affected,
york	york,
förstod	understood,
förts	brought,
kommunala	local,municipal,
tempererat	temperate,
tyst	quiet,
inleds	starts,
barns	childrens,
via	through,
area	area,
banor	paths,line,
david	david,
benämnas	named,
strida	fight,
krets	circuit,
helst	rather,
tvserier	tv shows,
nivå	level,
austin	austin,
revolutionens	the revolutions,
stämmer	correct,
isbn	isbn,
ursprungsbefolkningen	the native population,
brasilien	brazil,
uppger	states,
åring	year old,years,
jesus	jesus,
skyddade	protected,
nätverk	network,
värdefulla	valueable,
omständigheter	circumstances,
veckan	the week,
kantonerna	cantons,
meddelanden	messages,
upphört	ceased,
kulturarv	cultural heritage,
rösträtt	right to vote,
demonstrationer	demonstrations,
teatern	the theater,
valda	chosen,
viktor	viktor,
juli	july,
tätorter	conurbation,
hasch	hashish,
sjögren	sjögren,
styrelseskick	government,
framgångsrikt	successful,
släkten	the family,
dödligheten	mortality,
bevarats	protected,
definieras	defines,
franske	the french,
arbetade	worked,
birgitta	birgitta,
uteslutande	exclusivly,
framgång	success,
sakta	slowly,
osmanska	osmanian,
franskt	french,
mälaren	mälaren,
tyskarna	the germans,
vecka	week,
hänvisning	reference,
aristoteles	aristoteles,
fyrtio	forty,
cohen	cohen,
anpassat	adapted,
avgörs	decided,
basist	bassist,
mil	swedish miles,
lopp	race,
ansåg	thought,considered,
filosofin	philosophy,
skick	state,
benämning	term,name,
protesterade	protested,
linda	linda,
lån	loan,
konstverk	work of art,
centra	center,
konkurrerande	competing,
centre	centre,
runorna	the runes,
who	who,
kungliga	royal,
missionärer	missioners,
efternamn	lastname,
tyskar	germans,
republikanska	republican,
undersökte	investigated,
generna	the genes,
tidskrift	newspaper,
upphovsrätten	copyright,
moberg	moberg,
styrka	power,
utgångspunkt	starting point,
återfanns	was rediscovered,
inhemsk	native,
uppdelade	divided,
manchester	manchester,
planerat	planned,
parken	the park,
eiffeltornet	the eiffel tower,
järnvägen	railroad,
asterix	asterix,
östfronten	the east front,
rytmiska	rhythmic,
satan	satan,
gemensam	common,
härskare	ruler,
piano	piano,
allmänhet	general,
snitt	on average,
lägger	lies,
fotbollsspelare	football player,
inflytelserika	influential,
bonde	farmer,
klassiskt	classical,
presley	presley,
närstående	kindred,
mun	mouth,
britterna	the brits,
ingredienser	ingredients,
mohammed	mohammed,
iranska	iranian,
nazitysklands	nazi germany,
influensa	influenza,
debuterade	debuted,
vänt	turned,
universitetet	the university,
national	national,
priset	the prize,
förbinder	connects,
europa	europe,
bön	prayer,
hinner	have time to,
författarskap	the writer,authorship,
nationernas	the nations,
anlände	arrived,
wembley	wembley,
bör	should,
sjönk	sunk,
ken	ken,
balansen	the balance,
översikt	overview,
industrialisering	industrialization,
sovjetiska	soviet,sovjet,
hårdare	harder,
utformning	layout,
förklaringar	explanations,
jon	jon,
barrett	barett,
konservativa	conservative,
marknaden	the market,
återförening	reunion,
påtagligt	substantially,
la	la,
vulkaner	volcanos,
nyare	newer,
vattnets	the waters,
tillgången	access,
tätbefolkade	densely populated,
kommendör	commandor,
klasser	classes,
jersey	jersey,
torn	tower,
demens	dementia,
dör	dies,
malcolm	malcolm,
leipzig	liepzig,
befogenhet	warrant,
stabila	stable,
styrkor	strenghts,
publicerat	published,
liberala	liberal,
utkom	issued,
keltiska	celtic,
företaget	the company,
kopplade	connected,
beskrivning	description,
månar	moons,
reaktorn	reactor,
växt	plant,
genetik	genetics,
företagen	the companies,
ämbetsmän	bailies,
naturtillgångar	natural resources,
regelbundet	regularly,
pengar	money,
nickel	nickel,
västmakterna	western powers,
bär	carryng,berries,here,
strömningar	sentiments,
tillämpar	administers,
gärning	deed,
prestigefyllda	prestigious,
kanarieöarna	the canary islands,
godkännande	approval,
bråk	fights,
augusti	august,
officiell	official,
anpassa	adjust,
könsorganen	the reproductive organs,
fördelade	divided,
erhöll	recieved,
rikets	the realms,
demokrati	democracy,
avrättades	was executed,
reaktion	reaction,
aktivitet	activity,
ondskan	the evil,
förlopp	process,
gemensamt	in common,
syftar	refers,
rättigheter	rights,
flickor	girls,
måleri	painting,
partner	partner,
alfabetisk	alphabetical,
uppstå	develop,
parti	party,
friidrott	track and field,
varar	lasts,
buddhism	buddhism,
pojkar	boys,
terrorism	terrorism,
anka	anka,
material	material,
columbia	colombia,
sade	said,
införa	introduce,
nederlag	defeat,
anfield	anfield,
student	student,
sorter	kinds,
kallas	called,
representera	represent,
flickan	the girl,
grenar	branches,
spåren	the tracks,
väger	weighs,
ekosystem	ecosystem,
onda	evil,
störta	rush,
summan	the sum,
sänds	sends,
mystiska	mystical,
sofie	sofie,
flertal	majority group,
förtroende	confidence,
miljöer	environments,
antisemitism	antisemitism,
rocken	rock,
reformer	reforms,
hoppa	drop out,
landområden	land areas,
kontinuerligt	continous,
fyller	turns,
filmens	the film's,
dess	its,
vanligare	more common,
historia	history,
tillverkning	production,
historik	history,
klassificering	classification,
lika	alike,
dubai	dubai,
vulkaniska	vulcanic,volcanic,
budet	the bid,
vallhund	herding dog,
djupa	deep,
symptomen	the symptoms,
scientologikyrkan	church of scientology,
regeringar	governments,
säkra	safe,
starkaste	the strongest,
gäst	guest,
homo	homo,
export	export,
skorpan	crust,
högst	highest,
transport	transportation,
gammalt	old,
kaspiska	caspian,
operation	operation,
hyser	accomodates,
tänker	thinking,
stieg	stieg,
låten	the song,
sålt	sold,
sjunker	sinks,
äta	eat,
symbol	symbol,
viggo	viggo,
ställningar	positions,
samlades	collected,
uppvärmning	heating,warming,
ateist	atheist,
reza	reza,
svaga	weak,
slut	end,
biologi	biology,
sommarspelen	summer games,
svagt	weak,
beredd	prepared,
ljung	heather,
television	television,
låna	borrow,
upplöstes	dissolved,
användande	use,
nordkorea	north korea,
kontinenten	the continent,
freedom	frihet,
angeles	angeles,
troligen	likely,
alexanders	alexanders,
mytologi	mythology,
socken	parish,
omgiven	surrounded,
potatis	potato,
monarken	the monarch,
återvänt	returned,
någorlunda	fairly,
planetens	the planets,
tillbringade	spent,
kristus	christ,
floden	the river,
vidta	take,
ljusare	lighter,
framtiden	the future,
emi	emi,
hammarby	hammarby,
födelsetal	birth rate,
val	choice,
densamma	the same,
museum	museum,
upprättas	establish,
peters	peters,
skola	school,
pjäser	plays,
jah	jah,
föga	little,
förändrades	changed,
distinkt	distinctive,
klockan	clock,o'clock,
fru	wife,
brand	fire,
bröder	brothers,
neutral	neutral,
radioaktivt	radioactive,
bud	bid,
stadens	the citys,
utrymme	space,
volvo	volvo,
lissabon	lisbon,
stormakt	great power,
monument	monument,
inrättades	established,
innanför	inside,
minuter	minutes,
missnöjet	grievance,
kuriosa	trivia,
hästens	horses,
stormakter	world powers,
ordbok	dictionary,
utöva	exercise,
tolkningen	interpretetation,
omloppsbanor	orbits,
krav	requirement,
månader	months,
öga	eye,
illinois	illinois,
distinkta	distinct,
lutning	closing,incline,
book	book,
arbetskraft	labor,
befolkningstillväxten	the population growth,
picchu	picchu,
ljuset	the light,
effektiva	effective,
intresse	interest,
serbiska	serbian,
francisco	fransisco,
behandlas	treated,
fira	celebrate,
uttalade	spoke,
astronomi	astronomy,
klar	done,
förhandlingar	negotiations,
bröt	broke,
akademisk	academical,
stad	city,
upprepade	repeated,
stan	town,
hjärnan	the brain,
stam	tribe,
inspiration	inspiration,
syskon	siblings,
nödvändigtvis	necessarily,
svag	weak,
dave	dave,
praktisk	practical,
inser	realizes,
nederländska	dutch,
alkohol	alcohol,
blogg	blog,
