ödleblad	houttuynia
zirkon	zircon
foster	fetus
fritid	leisure
havskattfiskar	anarhichadidae
flicka	girl
makadam	macadam
befruktning	fertilisation
ängssyra	sorrel
ökenråttor	gerbil
neologi	neology
byrå	bureau
häcklöpning	hurdling
fröväxter	spermatophyte
rorsman	helmsman
brushane	ruff
högtryck	anticyclone
bläckpenna	quill
resurs	resource
eker	spoke
sugga	sow
mellanfot	metatarsus
koprolali	coprolalia
mullusfiskar	goatfish
metionin	methionine
långbåge	longbow
georgier	georgians
biogeografi	biogeography
depolarisering	depolarization
producent	producer
frekvens	frequency
stätta	stile
privilegium	privilege
akondroplasi	achondroplasia
besserwisser	know-it-all
promemoria	memorandum
fagocyt	phagocyte
geomorfologi	geomorphology
reologi	rheology
monografi	monograph
bioetik	bioethics
väska	bag
plattform	platform
kvast	broom
motorväg	autobahn
draperi	drapery
aktiv	active
gräslök	chives
azidgrupp	azide
stolpiller	suppository
ingenjör	engineer
laryngoskop	laryngoscope
kampanil	campanile
spindlingar	cortinarius
fåfotingar	pauropoda
klimatologi	climatology
fotbeklädnad	footwear
kupol	cupola
konsubstantiation	consubstantiation
giftsnokar	elapidae
baptism	baptist
nätvingar	neuroptera
schack	chess
sats	sentence
hällristning	petroglyph
kombattant	combatant
höftledsgrop	acetabulum
maffia	mafia
likör	liqueur
gom	palate
antropogen	anthropogenic
peang	hemostat
rubrik	rubric
reduktion	reduction
loggbok	logbook
rede	nest
