foster	,mrs. foster,infant,fomentar,fetuses,foster,do not need,nothing,embryonic,fetal
schack	schack,zircon,shack,performance,execution,check
loggbok	log book,analogue,log
stätta	,start,stood,allow,created
resurs	resusrs,resurs,factory,resources
monografi	every,thesis,each
koprolali	,number,coporolalia
mullusfiskar	,mullusfiskar (fish),mullets,don't know what it is except for a kind of fish,fish,mullusfiskar,admit,accept,mullisfiskar (fish),allow,red mullet,mullet,goatfishes
kvast	factories,groom
sugga	,coins,barrier,block
mellanfot	,metatarsals,mellanfot,metatarsel,islands
fagocyt	,fagocyt,phage,fagocyte,way
draperi	acoording,corresponding,drapery; curtain,curtains
reologi	,ether,reologi,air
fotbeklädnad	chaussure,shoewear,foot gear,chausurre,replacement
ökenråttor	,Ökenråttor,known,Ökenrättor,famous,gerbils; desert rats,ökenrättor
reduktion	processes
rubrik	title,many,header,quite a few,riburk,runrik,head line; rubric,heading
peang	,clamp,evolution,forceps,hemostatic clamp,hemostatic forceps,peang
azidgrupp	,azido group,lost,amide,azite group,azidgrupp
ödleblad	,Ödleblad,dleblad,lizard blade,houttuynia cordata,colour,lizardtail,odleblad,lizardleaf,ödleblad,color
sats	covering,theorem,cover,rate,proposition,statement,sets,proof,theorems; sets
befruktning	judaism,fertilizing,stimulation,conceptions,befrukning,conception,monograph
makadam	metal,trip,congress
flicka	pocket,jewish
fåfotingar	,over,centipede,n/a,arthropods,dafotingar,fÃ¥fotingar,fafotingar,pauropods
spindlingar	,slindlingar,cortinariuses,webcap,spindlingar,fungus,stalin,cortinarus,spiders,this is not a swedish word.
väska	,kazan,fluid,suitcase,vasks,its,pan
fritid	records,spare time,recreational,leisure time; spare time,record
bioetik	biotik,,bio ethics,wars,warrior
höftledsgrop	,hoftledsgrop,concave joint surface,mineral,hip pit,hip joint,aetabulum,hip joint fossa,minerals,ores
neologi	neologism,,plans,projected,neologi,planned,girl
långbåge	,long arc,i think it is language, but spelt incorrectly below.,many,ships,angbage
akondroplasi	,archondroplasia,created,achodroplasia
brushane	,secondary,rushane,brushane (bird)
antropogen	conference,man-made,anthropogeny,ntropogen
häcklöpning	,hackopning,hurdles race,hurdle,hacklopning,coin,hurdle-race
stolpiller	,web,pauropoda,network,suppositary
gom	related,corresponding,market organization,gum
frekvens	date,freckvens,by number of,value
geomorfologi	,stability,stable
ingenjör	complex,hard,ingenjor
producent	pregnancy,producers,produce,producent; tillverkare
depolarisering	depolarisation,,de-polarizing,nikolayevich,nikolaevich
maffia	,clinically,clinical,the mob
fröväxter	,about,provaxter,phanerogams,seedlings,spermatophytes,with
laryngoskop	,laryngoscopes,evolution,llaryngoscope
georgier	,the georgians,georgier,about, approximate
biogeografi	,evolution,use,usage,biogegraphy,biogeografi
likör	financing
privilegium	oh,privelege,privlege,privileium,privledge
rede	,clutch,ways,coated,means of
rorsman	,usage,rosman,helms man,using
motorväg	high way,tiumen,tyumen
metionin	,founded,creation,mentionin,created
högtryck	,high presssure,flat out,the heat is on,hotryck,high pressure,pressure,he
kupol	,regularly,combatant,regular,cu
kampanil	,kampanil,castle,lock,phagocyte
giftsnokar	,elapidaes,venomous conks,venomous grass snake,poison snakes,venomous snakes,elipidae,giftsnoakar,venomous snake,located,venom,passed,toxic snooping,venom snooping
zirkon	further,assisted,contributed
konsubstantiation	,no idea what it means,konsubstantiaion,korea,consubstantion,konsubstantiation,con-substantiation
hällristning	,halristning,chives,stone carving,agency,rock engraving,n/a,agencies,rock,rock engravings,venom snooping
ängssyra	,suppress,Ängssyra,sorell,suppression,sorrels,angssyra (perennial herb)
klimatologi	,use,klimatology,have,climateology
plattform	lost,platform; stand,platform, pad, stand,stage; platform,the plates,old plate,plattform
gräslök	chive,culture,raslok
besserwisser	,a,pundit,give,smartass,bewiseacre,exact: better knower; equivalent: know-it-all,between
nätvingar	,(nätvingar) an order in the class insects.,natvinger,lacewings,neuropteran,net wings, it's a animal,each,nätvingar,netwings,lacewing,natvingar
baptism	,universe,the universe,döpare
havskattfiskar	,catfishes,congress,havskattfskar,catfish fish,ocean catfish,seawolf,mullet,have duty fish
bläckpenna	statistics,ball point pen,ink pen,ink,ball point pen; pen,balck pen,black pen
promemoria	short essay,,aide-memoire,stalin,pm; memorandum,pormemoria,promemoria
