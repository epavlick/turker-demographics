vanligast	most,most usual,most common,
nordisk	nordic,
uppemot	almost,up,
stammarna	tribes,strains,
arternas	the species,species,
jihad	johad,jihad,
elva	eleven,
invandrare	immigrants,immigrant,
hållas	be,be held,
albumet	album,
slå	beat,hit,
albumen	the albums,albums,
hermann	hermann,
lord	lord,
vann	won,
lyckats	succeeded,
dela	divide,dividing,
katoliker	catholics,
syrgas	oxygen,
regional	regional,
upptar	occupies,
portugals	portugal,
dels	both,
skicklig	skillful,proficient,skilled; skillful,
statlig	state,government,
medelhavet	mediterranean sea,mediterranean,
andre	other,
helsingborg	helsingborg,
haber	haber,
befogenheter	authorities,powers,
triangelns	triangle,
flyr	flees,escapes,
urskilja	discern,
sovjetisk	soviet,
sture	sture,
sammansatta	composed,
ungerns	hungary,hungrarys,
hanar	males,
upprätthåller	maintains,maintaining,
åsikten	the opinion,view,
åsikter	opinions,
breddgraden	latitude,parallel,
fossil	fossil,
koffein	caffeine,caffein,
jönsson	jönsson,
filosofer	philosophers,
aten	athens,
hårda	hard,
biografi	biography,
vägrar	refuses,refuse,
filosofen	the philosopher,
motståndsrörelsen	the resistance,resistance,
regnskog	rain forest,rainforest,
baháulláh	bahaullah,bahullah,
föräldrarna	parents,
valrörelsen	election campaign,
bipolär	bipolar,
kids	kids,
demokratier	democracies,
naturen	the nature,nature,
blåser	blowing,
vicepresident	vice president,
robin	robin,
miljarder	billion,billions,
karin	karin,
systematiska	systematic,systematical,
unik	unique,
norsk	norwegian,
iis	ii's,
marino	marino,
hamas	hamas,
systematiskt	systematic,
ansluta	join,connect,
dna	dna,
sjukdomen	disease,
strikt	strict,
fuktiga	damp,damply,
betraktats	(been) viewed,
music	music,
dns	dns,
fuktigt	moist,damp,humid,
pjäs	piece,
musik	music,
befolkningstillväxten	the population growth,the growth of population,
mercurys	mercury's,mercurys,
holm	holm,
politiker	politicians,politician,
slutligen	back end,
bulgariska	bulgarian,
temperaturen	temperature,
kalksten	limestone,
rasen	the race,
teman	themes,
temperaturer	temperature,
ofta	usually,often,
avancerad	advanced,
vännen	the friend,friend,
köpa	buy,purchasing,
befolkningsutveckling	population development,population growth,
vågen	the wave,scale,
stommen	body,frame,the foundation,
köpt	purchased,bought,
passagerare	passengers,passenger,
kapitalismen	capitalism,
want	want,
absoluta	absolute,
vänner	friendas,friends,
igelkottar	hedgehogs,
hon	she,
kallare	colder,
hov	court,
how	how,
hot	hot,
pågick	lasted,
folkmusik	folk music,
typen	the type,type,
fylla	fill,
inrikes	domestic,
trettioåriga	13 year olds,
barbro	barbro,
sedd	seen,
objekt	object,
turkiet	turkey,turklet,
sankt	st.,sankt,
typer	characters,types,
stormaktstiden	great power period,greatness,
grekiska	greek,
isär	ice,apart,
arbeten	works,
deutsche	deutsche,
hemlandet	the home country,the homeland,
wind	wind,
skådespelerska	actress,
varv	revolutions,dockyard,
ormar	snakes,
vars	whose,
dalí	dali,
organismen	the organism,organism,
vare	either,
varg	wolf,
organismer	organism,organisms,
vara	be,
barnet	child,
mabel	mabel,
varm	hot,warm,
publicerade	published,
besläktade	related,
nutida	present(-day); contemporary,present,
wales	wales,
målade	painted,
assyriska	assyrian,
fil	master of,file,
avgå	resign,
väte	hydrogen,
hemlighet	secretly,darkness,
säljande	selling,
bestämmer	decide,
hänga	hang,
närliggande	adjacent,nearby,
silver	silver,
utvecklat	developed,evolved,
utlänningar	foreigners,
utvecklar	develops,development speaker,
utvecklas	development,
terrorister	terrorists,
tingslag	things type,
debut	debut,
utveckling	development,
tillgängligt	available,
utvecklad	developed,
andrew	andrew,
ingrid	ingrid,
tillgängliga	available,
uppnådde	met,achieved,
talade	spoke,
sapiens	sapiens,
angola	angola,
serier	comics,series,
allan	allan,
utvecklandet	development,
serien	the series,
truman	truman,
axelmakterna	axis,
varken	either,
kontrollerade	controlled,
slovenien	slovenia,
försökt	tried,
förändringar	changes,
foundation	foundation,
debatter	debates,
ian	ian,
anarkister	anarchists,
metallica	metallica,
arbetsplats	work,workplace,
ägnade	dedicated,
sannolikt	probably,probable,
att	that,
sysselsätter	employs,
atp	atp,
okända	unknown,
malmös	malmö's,malmö,
sydost	south east,southeast,
givetvis	course,naturally,
grannlandet	neighboring,the neighbouring country,
östberg	Östberg,ostberg,
tecknade	cartoon (-s),drew,
övre	upper,top,
djurgården	djurgården,zoo,
förespråkar	advocate,advocates,
xii	xii,
xis	the eleventh's,
master	masters,master,
vågade	dared,
ära	honor,glory,
bitter	bitter,
förändringarna	changes,change,
senaten	senate,
bokstäverna	the letters,letters,
förmögenhet	fortune,wealth,
placerade	placed,
nirvana	nirvana,
påverkad	influence,affected,influenced,
ahmed	ahmed,
skatter	taxes,
upphov	origin,source,rise,
tyckte	found,
påverkan	impact,influence,
tree	tree,
upplysningstiden	enlightenment,age of enlightenment,
nations	nation,nations,
påverkat	influenced,affected,
varje	each,
utformningen	the layout,
påverkas	affected,
tretton	thirteen,
obligatorisk	obligatory,mandatory,
folkmängden	population,
försörja	support,
densitet	density,
assistent	assistant,
kriterierna	criteria,
boston	boston,
dricker	drinking,drinks,
filosofisk	philosophical,philosophic,
halva	half,
joakim	joakim,
trakten	the region,region,area,
fasta	solid,firm; set; solid; fast; fasting,
kroatien	croatia,
krigsmakt	military power,armed forces,
östeuropa	eastern europe,east europe,
skaffa	obtain,gain,
förhärskande	prevailing,
hjälpmedel	aid,means agent,
bedrivs	conducted,
katalonien	catalonia,
konserthus	concert hall,concert,
victoria	victoria,
gallagher	gallagher,
medlemsstaterna	member states,
anteckningar	notes,
bedriva	carry,prosecute,
eftersom	because,
thriller	thriller,
övertog	took over,overtook,
annars	else,
singer	singer,
morgon	tomorrow,morning,
arkitektur	architecture,
öland	oland,öland,
camp	camp,
utmärkande	characteristic,distinguishing,
förlorar	loss,loses,
översatt	translated,
förlorat	lost,
grovt	heavy,rough,roughly,
passerade	passed,
singel	single,
tänkte	thought,was going to,
inspelning	recording,
ungar	kids,kids; offsprings; young,
representanter	representatives,
anorektiker	anorectics,anorexic,anorectic,
bandmedlemmar	band members,
konkret	specific,concrete,
pris	price,
teater	theatre; theater,theater,
louise	louis,louise,
populärkultur	popular culture,
buss	bus,
than	than,
övergår	surpasses,released,
sekulär	secular,
bush	bush,
omvända	reverse,
rice	rice,
mottog	received,
lastbilar	truck,
storbritanniens	united kingdom,
tillståndet	state,condition,the state,
rättegången	trial,the trial,
årsdag	anniversary,
metoder	methods,
upprätta	establish,up,
metoden	the method,
dansk	danish,
plats	place,place; position,
nathan	nathan,
lyssna	listening,listen,
begravning	funeral,
innebörd	meaning,
spänning	voltage,
hantverk	crafts,
×	x,
kallt	cold,coldly,
sköta	operate,handle,
utgåvan	the edition,
uppgift	task,data,
framfördes	framfordes,were,
kontroll	control,
release	release,
kalla	cold,
ovtjarka	caucasian shepherd dog,
blev	became,was,
etik	ethics,
flagga	flag,
skulle	could,would,
skriva	write,
bygger	based,
arlanda	arlanda,
skrivs	written,printed,
nuförtiden	nowadays,
hedersdoktor	honorary degree,honorary doctorate,
manson	manson,
förhindra	prevent,
wikipedia	wikipedia,
upphovsrätt	rise knob,copyright,
sundsvalls	sundsvall,(city of) sundsvall's,
figur	figure,
sista	last,
siste	last,
österrike	austria,
ringa	call,
rollen	role,the role,
henrik	henrik,
ställning	position,
lanserades	launched,was launched,
tilldelades	awarded,
kommunikation	communication,communications,
världsturné	world tour,
roller	roles,
yttre	outer,
tillämpar	practice,administers,
tillämpas	applied,
huvudet	head,the head,
country	country,
sparta	spartans,sparta,
följas	followed,
pitt	pitt,
edgar	edgar,
nordiska	nordic,
anordnas	provided,arranged,
nordiskt	nordic,
genus	gender,genus,
logik	logic,
summan	sum,the sum,
igelkotten	the hedgehog,
folkmordet	genocide,
armén	the army,
herr	mister,mr,
afrikanska	african,
fra	fra,
union	union,
avgörande	settling,decisive,essential,
fri	free,
tiotusentals	tens of thousands,
operationer	operations,
socialistiskt	socialistic,socialist,
årtionde	decade,
fru	mrs.,wife,
arbetslösheten	unemployment,
verktyg	tool,tools,
barndom	childhood,
life	life,
café	cafe,café,
huvudstäder	capitals,
ändrade	changed,modified,
arkiv	archives,archive,
närvarande	present (-ly),present,
dave	dave,
kometer	comets,
chile	chile,
övergripande	over arching,overall,general,
chili	chili,
parterna	parties,
intag	intake,
slutliga	evenutal,ultimate,
frankrikes	frances,
castro	castro,
klarade	passed,
organisera	organize,organizing,
kontraktet	the contract,contract,
tintin	tintin,
åke	åke,
brister	failures,inabilities,
gärna	i'd love to,readily,
desto	the,ever,
stämma	meeting,
player	player,
fascismen	the fascism,fascism,
australia	australia,
bristen	lack of,lack,
slag	kinds,type,
madonna	madonna,
tät	compact,sealed,frequent,
serbisk	serbian,
tillhandahåller	provides,
vrida	twist,turning,
foton	images,photos,
agnetha	agnetha,
european	european,
materiell	material,
funktionen	function,the function,
josef	joseph,josef,
topp	top,
värde	value,
emi	emi,
tunn	thin,
föras	be,be brought,taken to,
synder	sins,
tung	heavy,
obligatoriskt	mandatory,
finska	finnish,
lucas	lucas,
kampanj	campaign,
centraleuropa	central europe,
gudinnan	the godess,
grundlag	constitution,
försvarade	defended,
manteln	mantle,
snö	snow,
köra	run,drive,
koloniseringen	colonization,
capitol	capitol,
dödsoffer	casualty,death victim,
biskop	bishop,
krigsmakten	armed forces,
körs	driven,being driven,
birmingham	birmingham,
utrotning	extinction,extermination,
valutan	currency,
kommunal	communal,municipal,
döda	dead,
givit	gave,
matteus	matteus,
han	he,
grafit	graphite,
vetenskapsmän	scientist,scientists,
bnp	gdp,
ideal	ideals,
muhammeds	muhammad,muhammed's,
huvud	head,
hette	name was,named,
lunginflammation	pneumonia,
har	is,has,have,
hat	hatred,
hav	seas,sea,ocean,
präst	priest,
underliggande	underlying,
svensson	svensson,smith,
narkotika	drug,narcotics,
livsstil	life style,lifestyle,
dagar	says,day,days,
melodifestivalen	eurovision song contest,
uppmärksammade	observed,noted,
county	county,
bobby	bobby,
sedlar	bills,
alice	alice,
konsert	concert,
residensstad	city of residence,county seat,
sebastian	sebastian,
ola	ola,
old	old,
företräder	preferred trades,representing,
people	people,
reagera	reacting,reaching,
parlamentarisk	parliamentary,
delade	split,
kulmen	culmination,the acme,peak,
fot	foot,ft,
for	for,
varierande	variable,varied,varying,
fox	fox,
angränsande	adjoining,adjacent,
utser	appoints,
utses	is appointed,designated,appointed,
akademi	academy,
idéer	ideas,
myndigheter	authorities,agencies,
annan	another,
neptunus	neptunes,neptune,
stefan	stefan,
påminner	reminds,out,
hörde	heard,
binder	bind,
olympiska	olympic,
möjligheterna	possibilities,the possibilities,
myndigheten	the authority,authority,
annat	alia,other,other; another,
evangelierna	gospels,
army	army,
mynnar	opening,
stjärna	star,
misstänkt	accused,suspect,suspected of,
nixon	nixon,
tillverkare	manufacturer,
hänt	suspension,happened,
delvis	partial,partly,partially,
döpte	renamed,
psykiska	psychic,mental,
marshall	marshall,
som	as,which,
sol	sun,
lagliga	legal,lawful,
son	son,
psykiskt	psychic,mentally,
fci	fci,
delarna	parts,
artikeln	the article,
hantera	handle,
nova	nova,
säkerhetspolitik	safety policy,security,
joseph	joseph,
homo	homo,gay,
fria	free,
jane	jane,
 mm	millimeter,
happy	happy,
saltkråkan	salt crow,
jönköpings	jönköpings,
offer	victims,victim,
öppen	open,
förhållandet	the ratio,
förhållanden	relationships,conditions,
öppet	open,
verde	verde,
tigern	the tiger,
avsevärt	substantially,considerably,
förväntningar	expectations,
drabbat	affected,
gymnasiet	high school,gymnasium,
drabbar	affect,troubles,
polska	polish,
syften	purpose,
pest	plague,
syftet	purpose,
fansen	fans,
moderna	modern,
liberal	liberal,
föregångare	predecessor,precursor,
konung	king,
lunds	lund,lund's,
låtar	songs,
modernt	modern,
krävde	demanded,
ericsson	ericsson,
elektromagnetisk	electromagnetic,
huvudperson	main person; main character,protagonist,
dotter	daughter,
protester	protests,
wallenstein	wallenstein,
republik	republic,
roll	role,
olja	oil,
reggae	reggae,
avskaffades	was abolished,
bostadsområden	residential,housing,residential areas,
palme	palme,
blått	blue,
vintrarna	the winters,
modell	model,
rolling	rolling,
utbildade	educated,formed,
danske	danish,
aragorn	aragorn,
tävling	competition,
noga	carefully,
sällan	rare,
povel	povel,
laddade	charged,
perioden	period,
kategorifödda	category born,category: born,
förtjust	fond,delighted,
trettio	thirty,
herren	lord,the lord,
perioder	periods; episodes,period,
time	time,
erkända	acknowledged,recognized,
skatt	tax,
erkände	confession,acknowledged,
oss	center,us,
ost	cheese,
uppgifter	information,tasks,data,
stödjer	support,supports,
avalanche	avalanche,
uppgiften	the task,task,
atombomben	atomic bomb,the nuclear bomb,
stålgemenskapen	steel community,
inkomst	income,
behåller	retain,
machu	machu,
vet	know,
fängelset	prison,
intresserade	interested,
grön	green,
vem	who,
framställa	represent; depict; produce,the installation,
bosnien	bosnian,bosnia,
musikstilar	music genres,music,
individer	subjects,
choice	choice,
individen	the individual,individual,
framställs	is depicted,prepared,
skillnaderna	the differences,differences,
kusterna	coasts,
initiativ	initiative,
lägre	lower,
inhemska	native,
saab	saab,
oppositionen	opposition,
team	team,
uppskattningsvis	approximately,
årig	year old,minor,
jämnt	even,evenly,
nybildade	newly formed,
scen	scene,stage,
sjunka	decrease,descend,
firandet	celebrate,the celebration,
måne	moon,
greve	count,earl,
känd	known,unknown,famous,
elton	elton,
köp	purchase,
kör	run,
kunskapen	the knowledge,knowledge,
beskydd	conservation,
axel	axel,
bosatte	settled,
kön	gender,sex,
kunskaper	knowledge,
bosatta	residents,
kusten	the coast,coast,
katter	cats,cat,
berättelsen	story,the story,
provinserna	provinces,the provinces,
galileo	galileo,
vintertid	winter-time,winter,
kuster	coasts,
katten	the cat,
huvudsakliga	main,
studien	study,the study,
genomgående	consistently,through,pervading,
hälft	half,
landslag	national team,
studiet	study,the study,
studier	studies,
love	love,
engelske	english,
styrkan	strength; unit; force,
publicera	publish,
kommit	come,
presenterade	presented,
canis	canis,
sprids	spreading,spreads,
samlat	collected,gathered,
samlar	collect,
positiva	positive,
änglar	angels,
vuxna	adult,
sprida	spread,
judarna	jews,
positivt	positive,
samlag	intercourse,
effektiv	effective,
ställt	taken,put,set,
ställs	is,
dagars	day,days,
hår	hair,
tillträdde	took,
ställe	stalle,place,
hål	hal,
ställa	make,set,installation,
tabellen	table,table; list,
dålig	poor,
grönt	green,
straffet	penalty,
kunskap	knowledge,
gröna	green,
phoebe	phoebe,
påvisa	detection,show,
stigande	rising,up,
locka	attract,
missförstånd	misunderstanding,misunderstandings,
locke	locke,
släktskap	relationship,kinship,
inkluderade	included,
rädda	save,lot of,
porträtt	portraits,portrait,
utnyttjade	utilized,
drama	drama,
milda	mild,
årligen	annually,yearly,annual,
skikt	layers,layer,
svenskan	swedish,
storleken	size,
trigonometriska	trigonometric,
européer	europeans,
levande	live,
riksdagen	parliament,the parliament,
gigantiska	gigantic,giant,
kungens	king,the king's,
löpande	running,assembly,
svart	black,
nyligen	recently,
data	data,
epost	e-mail,email,
portugisiska	portuguese,
stress	stress,
natural	natural,
bergarter	rock types,minerals,rocks,
undervisning	teaching,education,
påstod	claimed,said,
ss	ss,
sr	sr,
sv	south west,
vikt	weight,
st	saint,
sk	so called,known,
so	so,
sm	swedish championship,
sa	said,
vika	fold,
se	see,
resulterar	resulting,result,
vintrar	winters,
resulterat	resulted,resulted in,
professorn	professor,the professor,
kong	kong,
antingen	either,
allvarligt	serious,severe,
clinton	clinton,
irländsk	ireland,
torg	square,
ingvar	ingvar,
dialekter	dialects,
utsätts	exposed,
jim	jim,
tilldelats	assigned,awarded,
begrepp	term,concept,
ersätts	replaced,
faderns	his father,the father's,
monopol	monopoly,
personlig	personal,
britter	britons,
hos	in; with,with,of,
änden	end,spirit,
öppnades	were opened,was opened,opened,
äldste	elders,eldest,
musiken	the music,music,
äldsta	oldest,
matcher	matches,games,
nation	nation,
records	records,
matchen	the game,match,
kategoripersoner	category of persons,
kantoner	cantons,
kravet	requirement,the demand,
musiker	musicians,
atmosfär	atmosphere,atmospheric,
lockar	curls,
förväxlas	confused,mistaken,
sidor	sides,
säga	say,
skivkontrakt	record deal,record contract,
dominerar	dominate,dominates,
domineras	dominated,
runstenar	runestones,
sägs	said,
dominerat	dominated,
födelsedag	birthday,
prisma	prism,
dynamiska	dynamic,
greker	greeks,
står	standing,star,
förstöra	destroy,ruin; destroy,
väljas	elected,choose,
hinduer	hindu,hindus,
krav	requirement,conditions,demands,
kött	meat,cones,
riktigt	real,
ockupationen	occupation,
sjuka	disease,sick,
avgör	decides,determines,
riktiga	real,
bränder	fires,
internet	internet,
roterar	rotates,
bla	blah,among others,
sfären	spheres,sphere,
garantera	ensure,guarantee,
vård	vard,healthcare,
våra	our,
singlar	singles,
sålde	sold,
bytt	changed,traded,switched,
byts	changed,replaced,
sålda	sold,salda,
väster	west,
vårt	each,
pilatus	pilatus,pilate,
dramaten	dramaten,
byte	bytes,
byta	change,trade,
föreställning	performance,
fyllt	filled,
pund	pound,
artister	artists,performers,
punk	punk rock,para,
flandern	flanders,
solna	solna,
artisten	the artist,artist,
gordon	gordon,
främst	foremost; primarily; chiefly,all,primarily,
givits	given,
självklart	course,
satte	put,
hård	diffcult,hard,
potter	pots,
one	one,
slutet	end,
tsunamier	tsunamis,
hårt	hard,
open	open,
ont	bad,
urin	urine,
city	city,
kraftigare	greater,more powerfully,
flytande	floating,
teologi	teology,theology,
skådespelarna	actors,
råolja	crude oil,
intill	beside,adjacent to,adjacent,
sjö	naval,lake,
nästa	next,
williams	williams,
animerade	animated,
vilka	who; which; that,who,which,
tillräckligt	sufficient,
dalar	valleys,
irakiska	iraqi,irakish,
tillräckliga	insufficient,sufficient,
svenskarna	the swedes,
yttersta	supreme,highly,
provins	province,
dygn	day,
fiskar	fishes,fish,
uppenbarelser	revelations,
berlinmuren	berlin wall,
kamprad	kamprad,
motståndarna	the opponents,opponents,
tankar	tank,thoughts,
sak	thing,matter; case,substance,
san	san,
sam	co,
generation	generation,
konsekvenser	consequences,
argument	arguments,argument,
församlingar	parishs,assemblies,
say	say,
känslan	feeling,the feeling,sense,
allen	allen,
turner	tournament,
staden	city,the city,
priserna	prices,the prices,
skickades	was sent,sent,
takt	rate,
general	general,
styrelsen	the board,board,
zoo	zoo,
jefferson	jefferson,
massa	mass,
övrigt	other,
förändringen	the change,change,
föder	gives birth,
muslimer	muslims,
finlands	finlands,
sekreterare	secretary,
tränare	coach,
mynt	coins,coin,
religionen	the religion,
betyda	mean,
religioner	religions,
forskningen	the science,research,
rådets	council,
kontroversiell	controversial,
driva	operate,run,
förändras	changes,
inledningen	the beginning,the introduction,
ursprung	origin,root,
fredspriset	nobel peace prize,peace price,peace prize,
rykte	reputation,
färdig	pre,done,
drivs	driven,run,
rött	cane,red,
olagligt	illegal,
axl	axl,
genomförts	out,
beckham	beckham,
vart	each,
ledd	led,
dimensioner	dimensions,
dahléns	dahlen,
sjöss	sea,
antalet	number,the number,
stärkte	strengthened,
slog	hit,
hockey	ice hockey,
caroline	caroline,
carolina	carolina,
beatles	beatles,
kategorimusik	category music,
återvänder	returns,atervander,
inlägg	post,
beatrice	beatrice,
egentliga	actual,
platta	flat,
undersöka	study,research,
rörande	concerning,
spetshundar	tip of dogs,
ländernas	the countries,countries,
artist	artist,
råd	council,
enighet	unity,
översättningen	translation,
roger	roger,
ljudet	noise,
varna	alerting,
sträcka	distance,
monark	monarch,
erbjöds	offered,
dagsläget	present situation,current situation,
översättning	translation,
spetsen	edge; top,tip,
brännvin	schnaps,aquavit,
snabbare	rapid,faster,
behovet	need,the need,
up	i[,up,
nederbörden	precipitation,the precipitation,
skärgård	archipelago,cutting garden,archipelagos,
talman	spokesperson,speaker,
ordspråk	proverbs,proverb,
enhetlig	single,uniform,
utgörs	consists of,is,
förvaltning	management,administration,
källa	source,
kritiserade	critisized,criticized,
begränsningar	limitations,limits,
upplever	experiencing,experience,
kontrakt	contract,
utgöra	compose,make up,
kilometer	kilometer,kilometers,
revolutionär	revolutionary,revolutions,
små	small,little, small,
gäller	of,grating,
amerikanskt	american,
anledningarna	reasons,the reasons,
screen	screen,
fynd	finding; finds,findings,
antika	ancient,
amerikanske	american,the american,
awards	awards,
inverkan	influence,
amerikanska	american,
mariette	mariette,
basisten	bassist,basist,the basist,
skönlitteratur	nonfiction,fiction,
mans	man's,
nationell	national,
rekord	record,
mani	mani,mania,
tillsätts	added,appoints,
långsammare	more slowly,slower,
upproret	the upprising,rebellion,
klimat	climate,
hamnade	landed,ended up,
anta	assume; adopt,adopting,
drogs	was pulled,was,
därtill	thereto,
teddy	teddy,
farfar	paternal grandfather,grandfather,
west	west,
airlines	airlines,
bolag	company,
luft	air,
cupen	the cup,cup,
lidit	sustained,suffered,
lånat	borrowed,
förr	sooner; past,sooner,before,
formen	the form,form,
formel	formula,
sångerska	songstress,singer,
regimer	regimens,regimes,
warhol	warhol,
tillåter	allow,
tillåtet	allowed,
pernilla	pernilla,
former	forms,
landskapen	landscapes,landscape,
samling	concentration,collection,
representativ	representative,
landskapet	landscape,
friska	healthy,fresh,healty,
situation	situation,position,
föregångaren	predecessor,
peruanska	peruvian,
ive	i've,
aston	överraska, undra,aston,
bror	brother,
ekonomi	economic,economy,
tillåtelse	permission,allowed,
blad	leaves,
beteckna	denote,
ohälsa	disorders,
världsbanken	world bank,
ståndpunkt	standpoint,position,
träffat	met,
wilhelm	wilhelm,
otto	otto,
träffas	reached,
oceanen	the ocean,ocean,
ekologi	ecology,
ludwig	lugwig,
nationalparker	national parks,
singapore	singapore,
sägas	is said,said,
lindgrens	lindgren's,lindgrens,
följer	resulting,
förkortning	abbreviation,
senator	senator,
dsmiv	dsm-iv,
personlighetsstörning	personality disorder,
måla	target,
tillfälle	occasion,time,
gestalter	figures,
avser	regard,refers to,
avses	regard,referred,
ifrågasatt	questioned,
eller	or,
iraks	iraq,
gudomliga	divine,
summer	sommar,
förluster	loss,losses,
bokförlaget	bokförlaget,publisher,
berättelse	tale,story,'s re,
rest	remain,residual,rest,
koncentration	concentration,
spårvagnar	trams,
psykologisk	psychological,
likheter	similarities,similarity,
resa	travel,
libyen	libya,
förlusten	loss; defeat,loss,
judarnas	jews,
kastar	throws,
heliga	saints,holy,holy; holy,
sprider	spreads out,spread,spreads,
helige	holy,
miljon	one million,million,
instrument	intrument,
körberg	körberg,
sänka	lower,
infördes	introduced,
unikt	unique,
heligt	holy,heligit,
störst	most,
snart	soon,once,
vinkel	angle,
dark	dark,
regim	regimen,regime,
unesco	unesco,
litteraturen	literature,
skadade	wounded,damaged,
stammar	strains,stutters,tribes,
statsreligion	state religion,
framsteg	progress,
tvserie	tv serial,
carl	carl,
tsunami	tsunami,
ekonomier	economies,
stupade	fallen,killed,
fossila	fossilized,fossil,
inter	inter,
intet	nothing,no,
jobbar	work,
nämnas	mentioned,include,
domkyrkan	cathedral,the cathedral,
ursprungsbefolkning	native population,indigenous,
ekman	ekman,
kännedom	known,knowledge,
närheten	near,
björn	bear,
föreslog	suggested,
institutionerna	institutions,
ddr	ddr,
än	yet,than,
exil	exile,
inkluderar	include,includes,
cannabis	cannabis,
varsin	opposite,
är	is,
atomkärnor	nuclei,nuclear particles,
ingående	input,enter into,
katolsk	catholic,
långstrump	longstocking,
jacksons	jackson's,jacksons,jackson,
nivån	level,
medlemsstater	member,member states,member-state,
stone	least,
organisationen	the organization,
ace	ace,
herrlandslag	men's national team,women's national teams,
vissa	some,
populationen	the population,population,
befinner	is,placed; situated; positioned; are,
digerdöden	black death,the black death,
populationer	populations,
lyssnade	listened,
organisationer	organizations,
industri	industry,industrial,
visst	specific,certain,
regissör	director,
berger	berger,
upplevelser	experiences,
ronden	round,
bryts	breaks,
nationalencyklopedin	national encyclopedia,the national encyclopedia,
image	image,
säkerhetsrådet	security,
partiet	the party,portion,
bryta	break,
partier	portions,parties,
lätt	easy,
bergen	mountain,
het	hot,up to date,
företag	company,companies,business,
kallats	called,
förintelsen	holocaust,the genocide,
philadelphia	philadelphia,
evangeliska	evangelical,
söker	seeks out,
hel	full,
hem	home,back,
hamnen	harbour,the harbour,
sover	sleep,
enorm	huge,enormous,
hänger	hanger,
hänvisning	reference,
project	project,
dagen	day,
complete	complete,
hells	hells,
bevarat	preserve,preserved,
bevaras	are protected,preserved,
mick	microphone,mike (microphone),
kontroverser	controversies,
språkliga	linguistic,
bevarad	kept,preserved,
åttonde	eighth,
rush	rush,
sällskap	company,groups,
jamaicas	jamaicas,jamaica's,
hexadecimalt	hexa-decimal,hex,
kvartsfinalen	quarter finals,quarterfinals,
utmed	along,
vinkeln	angle,the angle,
afrodite	aphrodite,afrodite,
förbundsstat	federal,federal state,
produkt	product,
puls	pulse,
krona	crown,
ac	ac,
ab	ab,
brodern	brother,
johnny	johnny,
redovisas	reported,shown,accounted for,
gustafs	gustafs,gustaf's,
am	am,
al	alder,
bronsåldern	bronze age,the bronze age,
as	as,
beordrade	commanded,ordered,
övernaturliga	over natural,
av	of,
håll	ways,hold,
väsentligt	substantially,relevant,
testamentet	testament,
vore	would,were,
federala	federal,
rökning	smoking,
innehåll	content,contents,
svårt	hard,difficult,
belönades	rewarded,awarded,
isolerad	isolation,
svåra	answering,difficult,
avslöjade	revealed,
såsom	such as,
gifta	marry,married,
värt	worth,
koppar	copper,
gifte	married,
medverkan	participation,
kvarstod	remained,
kategorisvenskspråkiga	category swedish-speaking,
terra	terra,
medverkat	participated,
medverkar	contributes,contribute,
terry	terry,
vanliga	regular,usual,
forntida	ancient,prehistoric,
kommunen	municipality,
skador	damage,
århundradena	centuries,
beteckning	label,
adam	adam,
omgivningen	surroundings,ambient,
decennierna	decades,
original	original,orignal,
renässans	renaissance,
känslor	feelings,
släppt	released,relinquished,
släpps	released,
elektron	electron,
halsen	throat,the throat,
anpassning	adjustment,
myntade	coined,
års	years,
släppa	release,
likartade	similiar,similar,
 kmh	km/h,
norr	north,
skogarna	the forests,forests,
number	number,
pojkvän	boyfriend,
ullevi	ullevi,
tv	tv,
romanen	novel,
nederbörd	rainfall,precipitation,
to	to,
mildare	milder,mild,
belägg	coating,evidence,
th	th,
nord	north,
te	tea,
sättas	turn,added,
ta	to,take,
avlägsna	remove,
använder	using,uses,
arvet	the inheritance,heritage,
telefonen	phone,the telephone,
strand	beach,
utländsk	foregin,foreign,
sant	true,
ensamma	alone,
djurarter	species of animals,animal species,species,
borrelia	borreliosis,
muslimska	muslim,
utsåg	declared,appointed,
sand	sandy,
siffrorna	figures,numbers,
områdets	the area's,area,
harry	harry,
sann	true,
språkbruk	language (use); parlance; phraseology,parlance,language,
förmedla	pass; express; mediate,pass,
döttrar	daughters,
samoa	samoa,
påståenden	claims,assertions,
synd	sin,
dödsstraff	death penalty,
utökade	expanded,increased,
vägnät	network,
pass	an,
givaren	donor,the giver,dealer,
syns	visible,
richard	richard,
stängt	closed,
delen	part,
soldater	soldiers,
islams	islams,islam's,
leif	leif,
gjorts	made,done,
hänsyn	light,consideration,
full	full,
gruppen	the group,group,
själen	the soul,
arkeologiska	archaeological,
grupper	groups,
legend	legend,
motstånd	resistance,opposition,
äventyr	adventures,
hindra	hinder,stop,
traditionella	traditional,conventional,
exklusiv	exclusive,
traditionellt	traditional,
social	social,
action	action,
oftare	more often,more,
varelser	creatures,
medlemskap	membership,
kommunistpartiet	communist party,the communist party,
vid	by,in,
ordinarie	permanent,regular,
vii	vii,
vin	wine,
young	small,
juridiskt	legally,judicial,
vis	vis,wise,
kuiperbältet	the kuiper belt,the cuyper belt,
vit	white,
spelaren	the player,
motsatsen	the opposite,opposite,
biskopen	bishop,the bishop,
mors	mother,
petroleum	oil,petroleum,
underordnade	subordinates,
pearl	pearl,
sitter	is,serve,sit,
presenterades	presented,
rhen	rhine,
dödligt	lethal,deadly,
mora	mora,
bevis	certificate,evidence,
mord	murder,
ragnar	ragnar,
uppskattad	estimated,
berättade	told,
uppskattas	is appreciated,estimated,
uppskattar	estimated,estimates,
schweiz	switzerland,
undergång	doom,destruction,
socialt	socially,social,
inträffade	occurred,happened,
medelklassen	middle class,
science	science,
monoteistiska	monotheistic,
klp	klp,
sociala	social,
morgan	morgan,
kapitalism	capitalism,
studenter	students,
läkaren	the doctor,physician,
samväldet	commonwealth,the commonwealth,
jakob	jakob,
säljas	is sold,sold,
nordvästra	northwest,north western,
skadliga	harmful,deleterious,
huvudstaden	capital,
mellersta	middle,the middle,
states	states,
stater	states,
spansk	spanish,
järnvägsnätet	railroad network,rail,
information	information,
vägnätet	road network,
hugo	hugo,
uppfattade	perceived,
ansetts	considered,regarded,regarded; viewed (as),
uppnått	met,achieved,
lejon	lion,
riksdagens	the parliament's,the parliaments,
retorik	rhetoric,
fortsättning	continuation,continued,
hustru	wife,
produktionen	production,the production,
referens	reference,
lanka	lanka,
köpte	bought,
barnens	childrens,
komplext	complex,
anklagade	accused,
pucken	the puck,
komplexa	complex,
utvidgning	enlargement; expansion,enlargement,
hållit	held,maintained,kept,
nationerna	the nations,nations,
blommor	flowers,
trade	esterified,
östblocket	cheese block,
scott	scott,
kvinnors	women,women's,
aktiviteter	activities,activity,
anställda	employed,
radion	radio,
vietnamkriget	the vietnam war,vietnam war,
känsla	feeling,sense,
alla	all,everyone,
högskola	college,
protestanter	protestants,
caesars	caesars,
miljön	environment,the environment,
termen	the term,term,
filip	filip,
termer	terms,
allt	all,
alls	all,
få	have; make; few,gain,fa,
van	van,
isaac	isaac,
konstruerade	constructed,
samhällets	society,of society,
berömda	famous,
inleda	initiate,
källan	source,kallan,
beräkna	calculate,
producerad	produced,
inledande	initial,
produceras	produced,
producerar	producing,
grekisk	greek,
producerat	produced,
introducerade	introduced,
producerade	produced,
olycka	accident,disaster,
intåg	advent,
budskap	message,
målning	painting,
graviditet	pregnancy,
blodet	the blood,blood,
denne	his,
denna	that,
härrör	derived,
enstaka	occasional,single,
england	england,
populärt	popular,popularly,
absolution	absolution,
sydöst	south east,southeast,
doser	dose,
populära	popular,
blues	blues,
förespråkade	advocated,
kretsen	the order,circuit,
finner	found,finds,
uppfördes	was constructed,built,
återkomst	return,
omröstningen	vote,
kopplad	connected to,connected,
garvey	garvey,
avgick	retired,
research	research,
norska	norwegian,
uppstått	resulting,arisen,
sammanfattning	summary,
besökte	visited,
kopplat	coupled; connected,connected,coupled,
hallucinationer	hallucinations,
highway	highway,
medel	middle,medium,
sparken	park,gets fired,fired,
alltmer	increasingly,more and more,
beethoven	beethoven,
stjärnor	stars,
poeter	poets,
driver	run,drive,
båda	both,
både	both,
kostade	cost,
ålands	Åland island's,aland,
kärnkraft	nuclear power,nuclear,
poeten	the poet,
teknologi	technology,
service	service,
turistmål	tourist attraction,
gatorna	the streets,streets,
samlas	together,
målningar	paintings,
skolan	school,
w	w,
nivåer	levels,
besök	visit,
uppenbarelse	apparition,
principen	the principal,principle,
bidragit	contributed,
relationer	relations,
foten	foot,
skiftande	shifting,
spekulationer	speculations,
såg	see,saw,
gemensamma	joint,common,
avel	breeding,
liknas	compared to,likened,
liknar	similar,
tove	tove,
wallander	wallander,
saint	saint,
sår	wound,
missade	failed,
besläktat	related,
läggas	laid,added,
chefen	head,commendant; commander,
tappade	lost,
zeus	zeus,
striderna	fighting,
zeppelin	zeppelin,
moder	mother,
svår	severe,difficult,
grace	grace,
obama	obama,
organiseras	organized,
återkom	return,returned,
organiserat	structured,
niklas	niklas,
koncentrerade	concentrated,
marknadsekonomi	market,market economy,
freud	freud,
organiserad	organised,organized,
nikolaj	nikolaj,nicholas,
ägg	eggs,
äga	be,aga,
väljer	select,elects,
inkluderas	include,is included,
statyn	the statue,statue,
generationen	generation,the generation,
förstörelse	destruction,
inkluderat	included,including,
ägt	taken,
generationer	generation,generations,
astronomin	astronomy,
visats	shown,demonstrated,
 au	au,
framåt	forward,forth,
varianten	version,variant,
norstedts	norstedt's,collins,
kongokinshasa	kong kinshasa,democratic republic of the congo,congo kinshasa,
varianter	variants,varieties,diversities,
vinterspelen	winter games,
arabisk	arabic,
edison	edison,
sydostasien	south east asia,southeast asia,
brooklyn	brooklyn,
plan	flat,level,
kombinationer	combinations,
arter	species,
utsattes	subjected,exposed,
cover	cover,
kanalen	the channel,channel,
kanaler	channels,
monarki	monarchy,
arten	species,
kombinationen	the combination,combination,
golf	golf,
gold	gold,
omfattade	included,
falska	false,
presidentens	president,the presidents,
detalj	detail,
karaktär	character,
falskt	false,
richmond	richmond,
framgångar	successes,success,
existensen	existence,
betydelser	values,meanings,
jämföra	compare,
befolkningstätheten	state of the population,
wayne	wayne,
betydelsen	the meaning,significance,
jämfört	compared to last,compared,
kontor	office,
karakteristiska	characteristic,
genomgick	underwent,
gratis	free,
evolutionen	evolution,the evolution,
tekniken	techinque,art,the technology,
tekniker	technician,
actress	actress,
utbildningen	education,
föll	fell,
erkännande	recognition,
victoriasjön	victoria lake,lake victoria,
tanken	the thought,idea,
ledare	conductors,leader,
cry	cry,
populärmusik	popular music,
byten	byte,
allmän	general,
river	tear,
sköt	shot,
någon	someone,anybody,
kriterier	criteria,
ses	be,
ser	sees,
koranen	the quran,
sex	six,
sed	sed,thirst,
psykologiska	psychological,
uppkomsten	onset,
lyckas	successful,succeed,
järnväg	railroad,rail,railway,
sen	then,since,
något	any,something,
sorters	kinds,kinds of,
institutet	institute,
församlingen	congregation,
trey	trey,
guinea	guinea,
neutralitet	neutral,
fission	fission,
kejsarens	emperor,the emperor's,emperors,
stärkelse	starch,
alqaida	al-qaida,al-qaeda,
rita	draw,drawing,
europe	europe,
europa	europe,european,
påverkar	affecting,
giftermål	marrige,marriage,
medveten	aware,
avvikelser	abnormalities,deviations,derivations,
medvetet	consciously,conscious,
möts	meets,meet,
fame	fame,
stadsdel	district,
demografiska	demographic,demographical,
forskare	researcher,scientists,
bästa	the best,best,
medicinering	medication,
förändring	change,
bäste	best,
messias	messiah,
stå	stand,
halmstads	straw city,
kopia	copy,
samma	the same,same,
transeuropeiska	transeuropean,
upprättades	was established,
krisen	crisis,the crisis,
kriser	crises,
church	church,
allierade	allied,allies,
decennium	decade,
sommaren	summer,
koalition	coalition,
mått	measurements,measurement,
väntade	expected; were waiting,waited,
tillväxt	growth,
potentiellt	potential,
kyrilliska	cyrillic,
upprättas	established,establish,
blod	blood,
pågår	(in) progress,underway,
föranledde	brought about,led,
beskrevs	was described,described,
skönhet	beauty,
östafrika	east africa,
fire	fire,
mind	mind,
taube	taube,
hovrätten	court of appeals,the court of appeal,
fritz	fritz,
uppleva	experience,
fritt	free,
föreningar	compounds,
systematik	systematic,
handling	act,
framträder	stand,appear,
projekt	project,
budget	budget,
feminism	feminism,
individerna	subjects,
bestående	comprising,lasting,
brottslighet	criminality,crime,
pressen	press,the pres,
föreställa	pretend; imagine,imagine,
arbete	work,work; labor,
vol	v,
von	von,
owen	owen,
motors	motor,
teoretisk	theoretical,
erkänna	recognize,
slöts	signed,
lokaler	facilities,place,
korruptionsindex	corruption perceptions index,corruption index,
arbeta	work,working,
kritiker	critics,
barney	barney,
gärning	deed,
möjlighet	oppertunity,possibility,
omvandlas	converted,
omvandlar	converts,
skalet	shell,the shell,
tillkom	hold back,resided,
barnen	children,
arméer	armies,
kritiken	criticism,the criticism,
laddning	charge,
kategoriavlidna	category deceased,
snarare	rather,
republiken	the republic of,the republic,
republiker	republics,
skapade	made,created,
debatten	the debate,
kring	on,around,
ledarskap	leadership,
fyra	four,
vargar	wolves,
euro	euro,
normala	normal,
normalt	normally,
person	person,
kelly	kelly,
johan	johan,
kontakter	contact,contacts,
finansiellt	financial,
sannolikhet	probability,
tunnelbana	subway,
stränder	beaches,
släppas	released,be released,
telegram	telegram,
stockholms	stockholm's,stockholm,
finansiella	financial,
kontakten	connector,the contact,
mandat	mandate,
fascistiska	fascist,fascistic,
rebecca	rebecca,
festivalen	festival,the festival,
symbolisk	nominal,symbolic,
nordväst	north west,
festivaler	festivals,
jönssonligan	jönssonligan,jonssonligan,
tomas	tomas,
hennes	her,
format	shaped,format,
turnéer	tours,
teologiska	theological,
melker	melker,
avvisar	reject,
skara	city in south-central sweden (uppland),crowd,
samarbete	co,
ivar	ivar,
västsahara	western sahara,
samarbeta	co,
da	da,
funnit	found,
skarp	sharp,crisp,
utlösa	trigger,
informationen	the information,
patrick	patrick,
ivan	ivan,
alexandra	alexandra,
ulrich	ulrich,
vojvodina	voyvodina,vojvodina,
lenin	lenin,
saknar	lacks,lack(-s),
saknas	missing,
användbar	useful,
utvecklades	developed,
avskaffade	abolished,absolished,
nåd	mercy,grace,
läste	read,
öka	oka,increasing,
brasilianska	brasilian,brazilian,
trafiken	traffic,the traffic,
turnerade	toured,
religion	religion,
riksförbundet	national association,
säger	said,says,claims; says,
be	be,
norra	north,northern,
ugandas	uganda,
västra	vastra,
bl	bl,
vagnar	carts,carriges,
bo	living,
bk	bk,
plocka	pick,
engelska	english,
bokstav	character,letter,
ordning	system,
santa	santa,
by	by,village,
källor	source,
ideologin	ideology,the ideology,
bosättningar	settlements,
patrik	patrik,
soldaterna	soldiers,the soldiers,
dagligen	day,daily,
gemenskaperna	communities,community,
aggressiv	aggressive,
arméerna	armeerna,armies,
stuart	stuart,
fungerande	functioning,effective,
för	of,to; for,for,
papper	paper,
texterna	text,
inte	not,
inta	taken,
colorado	colorado,
syret	the oxygen,oxygen,
hemingway	hemingway,
efterföljande	subsequent,
spridas	spread,disseminated,
kraven	the demands,requirements,
popsångare	popsinger,pop singer,
uppkallad	named,
orsaken	reason,cause,
förlaget	publisher,
seger	victory,
veckor	weeks,
kategorimusikgrupper	category of music groups,
dröja	take,
utbröt	erupted,broke out,
samerna	sami,
knuten	tied to,bound,knot,
fattigdom	poverty,
förbindelse	connection,
européerna	europeans,
poster	positions,post offices,
rörlighet	mobility,movement,
pastor	pastor,
begreppen	the concepts,terms,
begreppet	the term,term,concept,
posten	post,
atom	atomic,atom,
kritisk	critical,
line	line,
lovade	promised,
lina	lina,
dröm	dream,syndrome,
fader	father,
cia	cia,
ut	out; up,out,
dom	conviction,
drogmissbruk	drug abuse, substance abuse, drug addiction,drug,
eddie	eddie,
ur	out,
konventionella	conventional,
distrikt	district,
uk	uk,
protestantiska	protestant,
galaxer	galaxies,
testamente	testament,will,
professor	professor,
översvämningar	flooding,
nämner	mentions,
härstammar	derived,stems,
diverse	miscellaneous,
utbyggt	develpoed,built,
makedonska	macedonian,makedonish,
nationalism	nationalism,
inblandning	involvement,incorporation,
matematiken	mathematics,
händelsehorisonten	the event horizon,place else horizon,
räkna	count,
värld	world,
edwards	edwards,edward's,
são	sao,
skrivits	down,
innehåller	contains,
nordafrika	north africa,
innehållet	content,
matematiker	mathematician,
siffror	figures,numbers,
upplaga	edition,
individuella	individual,
besegra	defeat,
dominerades	was dominated,dominated,
radikala	radical,
djurgårdens	djurgården's,
lucia	lucia,
ägnar	spend time,spends time,
konstantinopel	constantinople,
riskerar	could,risks,
springsteen	springsteen,
radikalt	radically,
slås	is hit,slas,
alltså	therefore,really,
land	country,
passagerarna	passengers,the passengers,
uppträdande	performance,appearance,conduct,
symtom	symptoms,symptom,
age	do,age,
texten	text,the text,
sawyer	sawyer,
texter	texts,
majs	corn,
förväntas	expected,
persbrandt	persbrandt,
släpptes	released,was released,
alltför	all too,way too,exessive,
bakåt	backwards,reverse,
turkisk	turkish,
dyraste	most expensive,
hamnar	lands,ports,
hamnat	ended up,got in to,
listade	listed,
dickinson	dickinson,
dancehall	dance hall,dancehall,
sent	late,
garden	garden,
märken	sign,
kedjan	chain,the chain,
palestinier	palestinians,
kommunistiska	communistic,communist,
flöde	feed,
drogen	the drug,drug,
känner	knows,
överleva	survival,
tillhörande	associated,belonging to,
magic	magic,
tro	believing,
påverka	impact,influence,
harbor	harbor,
eva	eva,
tre	three,
jobbet	work,the job,
romerska	roman,
överlevt	survived,
romerske	roman,
opinionen	opinion,
innebörden	meaning,the significance,
leonardo	leonardo,
bolsjevikerna	bolsheviks,the bolsheviks,
natur	nature,
regelbundna	regular,
ställde	set,stood up,asked,
årtionden	decades,
video	video,
förhållandevis	relatively,
legitimitet	legitimacy,
victor	victor,
antog	adopted,
index	index,
expressen	expressen,
anton	anton,
praktiken	effectively,practically,
indiens	india's,indias,
suveräna	terrific,sovereign,
möjliggör	enables,enable,
birk	brik,birk,
indian	indian,
ledande	conductive,leading,
wembley	wembley,
stadskärna	city core, city center,town,
led	suffered,step,
lee	lee,
lyckades	managed,succeeded,
upphovsrätten	copyright,
sålunda	thus,
leo	leo,
let	cleanly,
lev	lev,
hälsa	health,
talang	talent,
begravd	buried,
motorvägarna	highways,the highways,
tegel	brick,
casino	casino,
titanic	titanic,
förutsätter	assume,requires,assumes,
högste	supreme,highest,
insulin	insulin,
högsta	highest,
opinion	opinion,
sekel	centuries,
huvudvärk	headache,
emot	vis,
förlora	lose,
oxenstierna	the oxenstierna,oxenstierna,
mening	meanings,sentence,
indianerna	the indians,indians,
anatolien	anatolia,
andreas	andreas,
varmare	heater,warmer,
rico	rico,
illegal	illicit,
hemlig	secret,
elever	students,
godkänna	approve,
klaviatur	keyboard,
orkester	orchestra,
projektet	project,
existerade	existed,
författning	constitution,
samspel	teamwork,
ytterst	very; extremely,highly,
överlevande	survivors,survivor; survivors; surviving,
villor	villas,
edwall	edwall,
lokalt	locally,local,
bidraget	grant,
advokat	bar,
ortodoxa	orthodox,
lokala	local,
peka	point (at; to; in),point,
gustafsson	gustafsson,
upprätthålla	keep up,maintaining,
process	process,
artiklar	items,
etta	number one,first,one,
tryckta	printed,
high	high,
syre	oxygen,
hercegovina	herzegovina,
sydöstra	south east,
föregående	preceeding; previous,
halmstad	halmstad,
frågor	questions,
saknade	missed,missing,
delad	shared,divided,
övergrepp	assault,abuse,assult (-s),
latinska	latin,
hormoner	hormones,
delas	shared,divided,
delar	proportions,parts,
delat	shared,divided,
sydvästra	southwest,southwestern,
kriminella	criminal,
gunwer	gunwer,
amerika	american,america,
djurens	the animals,animal,
profeten	prophet,the prophet,
insatser	action,
regeringsmakten	govermental power,government power,
platt	plate,
väckt	brought,awaken,
slutsatser	conclusions,
gitarr	guitar,guitarr,
element	elements,
lundgren	lundgren,
nancy	nancy,
kvinnliga	female,
byggnadsverk	building,edifice,
borde	should,
handboll	handball,
diskar	disks,
houston	houston,
möjligt	possible,
hårdast	hardest,the hardest,
universiteten	universities,the universities,
frånvaro	absent,absence,
hunnit	had time to,
universitetet	the university,university,
bensin	gasoline,
sydligaste	southernmost,most southern,
möjliga	possible,
solvinden	the solar wind,solar wind,
västerbottens	västerbottens,west bothnia,
eliten	the elite,elite,
uppdelat	divided,split,
fristående	independent,stand-alone,
tecknet	the sign,sign,
uppdelad	divided,split,
puerto	puerto,port,
beståndsdelar	constituents,elements,
ovanlig	unusual,rare,uncommon,
konkurs	bankruptcy,
bekant	known,acquaintance,
bryter	breaks,breaking; violating,
hemmaplan	home,home turf; domestic (level),
dock	nevertheless,however,
utgår	deleted,
rotation	rotation,
huvuddelen	bulk,main part,
sönder	broken,probes,
peking	beijing,peking,
välfärd	wealth,welfare,
intressen	interests,
fortsätta	remain,continue,
smallwood	smallwood,
fördrevs	was banished,ford described,
burton	burton,
books	books,
intresset	the interest,
frac	fraction,
bay	bay,
etymologi	etymology,
matrix	matrix,
borderline	borderline,
billiga	cheap,
utbildad	educated,
enskilda	individual,
anledningen	reason,therefore,
umgänge	intercourse,
kapitalismens	capitalism's,capitalism,
marxistiska	marxist,
bekräftades	was confirmed,
fram	until,out,
undertecknades	signed,
legat	formed,
redskap	device,tool,
egenskaperna	the qualities,properties,
mötte	motte,met,
sköts	postponed; run,shot,
påverkats	affected,
melankoli	melancholy,
uppe	up,(on) top, up, above,
förts	brought,cont,
tempererat	temperate,
dubbel	double,
liggande	placed,overhead,
kompositör	composer,
krävt	required,
våldsam	violent,
krävs	needs,requires,
david	david,
blanda	mix,
profeter	prophets,profets,
krets	sphere,circuit,
helst	rather,anyone,
hussein	hussein,
kräva	require,demand,
skillnad	difference,unlike,
playstation	playstation,
åring	year old,years,
komplicerade	complex,
jesus	jesus,
användningsområden	possible use,applications,
schweiziska	swiss,
muhammad	muhammad,
nordkoreanska	north korean,
studerade	studied,
värdefulla	valueable,value,
festival	festival,
system	system,
bygget	construction,
vänster	left,
hebreiska	hebrew,
tränga	permeate,cut in,
teatern	the theater,theater,
blivit	become,was,
utbyggnad	development,expansion,
havet	sea,
pristagare	laureate,
konservativ	conservative,
utländska	foreign,
haven	the seas,
visdom	wisdom,
hampa	hemp,
samverkar	co,co-operating,
roberto	roberto,
stewie	stewie,
roberts	roberts,
reagans	reagan's,reagan,
troende	believers,faithful,
vecka	week,
jonatan	jonatan,
räcker	enough,sufficient,
användaren	the user,user,
producent	producer,
förslag	'proposal,proposed,
flygplats	airport,
kritiskt	critical,
instruktioner	instructions,
mills	mills,
filosofin	philosophy,the philosophy,
sinatra	sinatra,
kritiska	critical,
best	best,
uppträdde	appeared,perform,occurred,
viss	certain,some,
finsk	finnish,
slutsatsen	concluded,the conclusion,
säkert	securely,
när	when,
nät	web,
trosbekännelsen	creed,
detta	that,
vardagen	the weekday,everyday life,
napoleons	napoleon,napoleon's,
visa	see,
uppror	rebellion,
flyga	fly,
förutsättningarna	prerequisites,conditions,
medan	while,
framgår	will be seen,is shown,
synliga	visible,
våren	spring,the spring,
bred	broad,
bokstaven	the letter,character,
face	face,
synligt	seen,
befolkningens	population's,population,
närmade	approached,
brev	letter,
beteende	behaviour,behavior,
uppdelade	divided,
manchester	manchester,
tyvärr	unfortunately,
hopp	hopes,hope,
fursten	prince,
östfronten	eastern front,the east front,
samisk	sami,
jan	jan,
simmons	simmons,
religionens	religion,religion's,
liksom	and,
jah	jah,
jag	i,
skarsgård	cut farm,skarsgård,
ilska	anger,
handla	act; buy; consume,act,
abba	abba,
parlamentet	the parlament,parliament,
lägger	put,lies,
fotbollsspelare	football player,footballers,
lucky	lucky,
generalen	the general,general,
bonde	farmer,
parlamenten	parliaments,
meter	meters,meter,
tidigaste	earliest,
britterna	the brits,british,
h	h,
rowling	rowling,
effekterna	the effects,effects,
iranska	iranian,
rymmer	has,holds,
guvernör	governor,
myndigheterna	authorities,the authorities,the authoroties,
debuterade	debut,debuted,
michail	michail,
konungarike	kingdom,
avlidit	died,
priset	the prize,rate,
kronisk	chronic,
lämplig	suitable,
freddy	freddy,
vietnams	vietnam's,vietnam,
författarskap	the writer,authorship,
sjöng	sang,
upprättandet	establishment,establishing,
längst	at,farthest,longest,
sjönk	sunk,sank,decreased,
balansen	balance,the balance,
värre	worse,
kategorisvenskar	category swedes,
striden	battle,fight,
finalen	final,
bolivias	bolivia,bolivia's,
strider	conflict,battles,
bilar	car,cars,
ende	only,
förklaringar	explanations,
kedjor	chains,
islamiska	islamic,
ett	a,one; a; an,
marknaden	the market,market,
figuren	the character,figure,
religiöst	religious,
beläget	located,base,
fåglar	birds,
egypten	egypt,
norge	norway,
etc	etc.,
marknader	markets,
ogillade	disliked,
belägen	situated,disposed,
utövade	exerted,exercised,
tätbefolkade	densely populated,populated,
ekvatorn	equator,the equator,
religiösa	religious,
framgången	success,the success,
co	co,
dör	dies,
ca	cirka,approximately,
mengele	mengele,
cd	cd,
död	dead,dod,
bröllop	brollop,
stabila	stable,
musikvideo	music video,
cp	cp,
öst	east,
dök	appeared,dove,turned,
antal	number of,number,
jussi	jussi,
keltiska	celtic,
företaget	the company,
moraliskt	morally,moral,
överallt	in all,everywhere,overall; everywhere,
kombination	combination,
rockband	rock band,
genetik	genetics,
moraliska	moral,
företagen	the companies,taken present,
antas	assumed,
antar	adopting,
typisk	typical,
frågorna	questions; issues,
molekyler	molecules,
tvungna	forced,forced to,
sänts	sent,
atlanta	atlanta,
haile	haile,
mandatperiod	term (of office),term of office,
långsamma	slow,
tjorven	tjorven,
rikets	its,the realms,
demokrati	democracy,
aktivitet	activity,
vd	ceo,
ondskan	the evil,
förlopp	process,developments,
omnämns	mentioned,is mentioned,
vi	we,
ryssland	russia,
vm	world championship,vm,
lust	desire,loss,
vs	vs,
flickor	girls,
skapare	creator,
föreligger	is,exist,
sitt	its,
slovenska	slovenian,
evenemang	event,
spela	play,
tupac	tupac,
armé	poor,
känt	known,
juan	juan,
medeltida	medival,medieval,
foundationthe	the foundation,
huden	skin,
paulo	paulo,
matthew	matthew,
und	und,
terrorism	terrorism,
flesta	most,
ball	ball,
columbia	columbia,colombia,
sade	said,
konstantin	constantine,
framförde	performed,presented,
nederlag	defeat,
anfield	anfield,
ikea	ikea,
sjukhus	hospital,hospitals,
diabetes	diabetes,
representera	represents,represent,
obamas	obama,obama's,
mänskligt	human,
klubbarna	the clubs,
väger	weighs,weight,
vägen	the road,road,
ledde	resulted,led,
ledda	led,
uno	uno,
versaillesfreden	versailles peace,treaty of versailles,
vägarna	paths,roads (roadways),
gatan	the street,
kontakt	plug,
paus	pause,paus,
aktuell	current,
renässansen	the renaissance,renaissance,
paul	paul,
pappa	dad,
tolkade	interpreted,
förknippas	associated to,
kunder	customer,
planeter	planets,
frågan	issue,the question,
englands	england's,
planeten	planet,the planet,
kosovos	kosovo,
filmens	the film's,
framtid	future,
förknippad	associated,
motorvägen	motorway,highway,
government	government,
ledarna	the leaders,conductors,
gul	yellow,
dess	then,its,
arbetarklassen	working class,the working class,
tillverkning	production,
pressas	pressed,
följeslagare	companions,companion,
lät	had,
emma	emaa,emma,
lär	teach,learn,
aktiebolag	companies,limited company; joint-stock company,stock company,
vallhund	herding dog,herder,
stadsbild	cityscape,
amazonas	the amazon rainforest,amazon,
symptomen	symptoms,the symptoms,
högskolan	hogs school,university,college,
flotta	fleet,
län	state,between,
tackade	thanked,said/thanked,
bredare	broad,
miniatyr|	miniature,
filmografi	filmography,
anarkismen	the anarkism,anarchism,
trotskij	trotskij,trotsky,
lägsta	lowest,minimum,
stannar	stop,stays,
transport	carriage,transportation,
skriftliga	written,
ockupation	occupation,
februari	february,februari,
kolonin	colony,
behandlades	treated,
flitigt	actively,frequent,
sålt	sold,
dags	time,
naturlig	natural,
kollektivtrafik	public transport,
ateist	atheist,
svaga	weak,
fråga	fraga,question,
förklaringen	the explanation,statement,
biologi	biology,
ateism	atheism,
östberlin	east berlin,
svagt	weak,
gandalf	gandalf,
smärta	pain,
vargen	the wolf,
användande	use,use; usage,
kontinenten	the continent,
må	mon,
erövrade	conquered,
höger	right,
blodiga	blooded,bloody,
angeles	angeles,
kontinenter	continents,
warner	warner,
solsystemets	solar system,
hittills	date,
burma	burma,
släpper	release,releases,
upplösningen	dissolution,disbandment,
sekelskiftet	turn,
planetens	planet,the planets,
kristus	christ,
lund	grove,
mera	more,
varma	hot,warm,
peters	peters,
skola	school,
blå	blue,blah,
fläckar	stain,
bedöms	expected,judged,
överbefälhavare	commander-in-chief,supreme commander,
tina	defrost,thaw,
radioaktiva	radioactive,
samlingar	collection,
förre	pre,
uppvisade	showed,
apollo	apollo,
radioaktivt	radioactive,
svält	starvation,starvations,
återkommer	will return,returning,
society	society,
official	official,
volvo	volvo,
ruset	the fuddle,intoxication,
stormakt	great power,
monument	monument,monuments,
inrättades	established,were implemented,
distribution	distribution,
ovanför	above the,above,
leukemi	leukemia,
heter	units,is named,
guy	guy,
utnyttjar	using,uses,
utnyttjas	utilized,used,
skilsmässa	divorce,
separerade	separated,
broder	brother,
banan	banana,
vitryssland	belarus,
månader	months,
sharia	sharia,
öga	eye,
distinkta	distinct,
särskilt	in particular,especially,
relationen	the relation,ratio,
månaden	the month,months,month,
modernistiska	modernistic,modernist,
bröd	bread,
övergång	transition,
francisco	fransisco,
uttalade	commented; made a comment; spoke about,spoke,
tider	times; ages,times,
förhandlingar	negotiations,
bröt	brot,broke,
tiden	time,
inspiration	inspiration,
syskon	sibling,siblings,
mozart	mozart,
sänker	lowers,lower,sinks,
tredje	third,
jordbävning	earthquake,
provinser	provinces,
kommersiell	commercial,
nederländska	netherlands,dutch,
brevet	the letter,letter,
näsan	the nose,nose,
child	child,
elisabeth	elisabeth,
bob	bob,
bosniska	bosnian,
tätort	urban,conurbation,
invadera	invade,
preussen	prussia,
konsekvenserna	impact,consequensis,
smålands	smaland's,småland,
bäst	best,
atlanten	the atlantic ocean,
bibel	insulin,bilble,
spel	game,
edward	edward,
grundande	founding,
ren	clean,
konsekvens	impact,consequence,
mördade	murdered,
konsekvent	consistent,consistency,
grönsaker	vegetables,
golvet	the floor,floor,
främsta	primary; foremost; primarily; principally,request,
främste	chief,premier,
geologi	geology,
jacob	jacob,
skolor	schools,
innefattar	comprises,includes,
uttryck	expression,
upphörde	ceased,
estland	estland,estonia,
jamaica	jamaica,
starkast	strongest,
ständerna	the cities,
galax	galaxy,
horn	horns,horn,
colorblack	color black,
alltsedan	since,
förbättringar	improvements,improvement,
eurovision	eurovision,
bakgrunden	background,
vidsträckta	broad,wide; broad,
kraftfull	forceful,
tolv	twelve,
bidrag	contribution,contributions,
vampyr	vampire,
cyklar	bicycles,cycles,
bidrar	contributes,
petra	petra,
musikalen	the musical,
räddar	saves,saved,rescues,
bortgång	passing,death,
pluto	pluto,
rapporterar	reports,
norstedt	norstedt,
begått	committed,
olsson	olsson,
studeras	studied,is studied,
sidan	page,side,
interstellära	interstellar,
regerande	reigning,ruling,
hänvisade	referred,
förblir	remains,remain,
stoft	dust,
träda	esterified,emerge,fallow,
placerades	placed,
akc	akc,
underverk	wonders,wonder,
kongressen	congress,
järnmalm	iron ore,
fastställdes	confirmed,set,
bro	bridge,
läkemedelsverket	medicines work,food and drug administration,
tillsammans	together,
faktiska	actual,
total	total,
bra	good,
stått	stood,
sarah	sarah,
ätten	the dynasty,dynasty,
negativa	negative,
foster	fetus,fetal,
indiana	indiana,
negativt	negative,
supportrar	supporters,
ifall	if,
förebyggande	preventive,
giovanni	giovanni,
fingrar	fingers,
award	award,
riksväg	national highway,highway,
nku	nku,
alces	alces,
inleds	starts,start,
kurderna	kurdish,kurds,
springer	running,
absorberas	absorbed,
friheten	freedom; liberty,freedom,liberty,
beväpnade	armed,
tänkare	thinker,
dokument	documents,
era	yours,era,
transparency	transparency,
specialiserade	specialized,special,
klorofyll	chlorophyll,cholophyll,
vietnamesiska	vietnamese,
gloria	gloria,
vackra	beautiful,fine,
felaktiga	false,
ekonomiskt	economic,economically,economical,
sommar	summer,
indien	india,
felaktigt	erronenous,error,
indier	indians,
enhet	unit,entity,
valborg	may day,valborg,
utlandet	abroad,
gotlands	gotland's,gotland,
solen	sol,
firas	celebrated,celebrate,
firar	celebrates,celebrate,
gillar	like,enjoy; like,likes,
leonard	leonard,
halland	halland,
beach	beach,
sammansatt	composed,compound,
rädd	scared,
biografer	movie theaters,movie theaters; cinemas,
kategorieuropas	category europe,
lag	law,act,
koreakriget	korean war,the korean war,
visste	did,
tjäna	profit,earn,make,
biografen	movie theater,cinema,
law	law,
orden	the words,words,
medlemsstat	member state,
vänsterpartiet	leftist party,left wing party,
lämningar	remnants,
green	green,
massmedia	media,
livets	life,life's,
ordet	word,
order	order,
arbetslöshet	unemployment,unemplyment,
natten	overnight,
office	office,
sovjet	soviet,
diagnos	diagnostics,
exempel	example,for example; for instance; sample(-s),
ramadan	ramadan,
söderut	south,
blandning	mix,mixture,
japan	japan,
bidra	contribute,
straff	punishments,
lagets	substrate,the team's,
fragment	fragments,
vanligtvis	usually,generally,
ämne	substance,
band	band,tape,
fredsbevarande	peace,peacekeeping,
bana	course,web,
they	they,
spelningen	the gig,
bank	bank,
ansvariga	charge,
huvudartikel	main article,
helvetet	hell,
dåliga	poor,bad,
diskuteras	discussed,
knutpunkt	hub,
tendens	tendency,
dåligt	poor,
område	area,
carlos	carlos,
erbjöd	offered,
germanska	germanic,germanian,
inflytandet	the influence,influence,
koldioxid	carbon dioxide,co,
voddler	voddler,
däggdjur	mammalian,
rummet	room,
kejserliga	imperially,imperial,
asteroidbältet	asteroid belt,the asteroid belt,
daniel	daniel,
därav	thereof,
trafik	traffic,
bruttonationalprodukt	gross national product,bnp,
oskar	oskar,
vete	wheat,
klimatet	environment,climate,
veta	know,out,
sedermera	subsequently,since,
veto	veto,
standard	standard,
förmodligen	probably,
tillbaka	back,
berör	affecting,affect,concerns,
amadeus	amadeus,
ange	set,
sprit	alcohol,
väldiga	immense,mighty,vast,
förefaller	appears,
professionell	professional,
väldigt	very,
höll	hold,gave,
personerna	people; persons,subjects,
funktioner	functions,features,
önskar	desired,desiring to,wish,
önskan	desired,
another	another,
statskupp	coup,
ingmar	ingmar,
synnerligen	remarkably; particularly,
drabbade	suffering,affected,
begränsas	limited,
begränsar	limit,limits,
ingen	no,
begränsat	limited,restricted,
sång	song,
lidande	sufferer,
växthusgaser	vaxthusgaser,greenhouse gas,
inget	not,no,
john	john,
begränsad	restricted,limited,
medborgare	citizens,
antisemitismen	anti-semitism,
äter	eat,eats,
varifrån	from where; wherefrom,from which,
albert	albert,
åland	Åland,
kvarvarande	lasting,remaining,residual,
persson	persson,
bojkott	boycott,
kraftverk	plant,power plant,
trupp	troops,troop,
zeeland	zealand,zeeland,
militära	military,
nedan	below,
symboliserar	symbolizes,
binda	tying,bond,
kronan	kronan,
sonen	the son,
scener	scenes,
används	use,
scenen	stage,
binds	bind,bound,
iron	iron,
byggts	built,
minut	minute,
använde	used,
använda	using,
årens	the year's,years,
skolorna	schools,the schools,
mannen	art,the man,
noterade	note,noted,
onani	masturbation,
höja	hoja,raise,
fåglarna	birds,
omvandling	transformation,
avancerade	advanced,
koloniala	colonial,
anledningar	reasons,
kalendern	calendar,calender,
stavning	spelling,
magnus	magnus,
höjd	height; above,height,
sjukvård	health care,healthcare,
aftonbladet	aftonbladet,newsweek,
lades	put,
figurerna	figures,characters,
närvaro	attendance,presence,
verkat	worked,acted,seemed,
verkar	acting,seems,
maiden	maiden,
bruce	bruce,
utställning	display,exhibition,
skansen	forecastle,
fjädrar	spring,feathers,
verkan	effect,
flygplatsen	airport,the airport,
aminosyra	amino acid,
vägg	wall,
eviga	eternal,
ägda	owned,
freja	joe,
ägde	tookplace; occured,was,owned,
bortom	beyond,beyond the,
läran	teaching,the teaching,
evigt	forever,eternal,
misslyckade	failed,
förväxla	confuse,mistake,
effekten	the effect,effect,
mitten	middle,
damer	ladies,
lewis	lewis,
hinduiska	hindu,
vanligen	usually,typically,
tilläts	was allowed,
effekter	effects; repercussions,effects,
fortplantning	reproduction,
vätet	hydrogen,the hydrogen,
sättet	manner,the way,
 kilometer	kilometer,
sätter	place,puts,sets,
näring	nutrition,
estetiska	aesthetic,
ambassad	embassy,
kejsar	emperor,
inställning	attitude,setting,
målvakt	goalee,goalkeeper,
variera	vary,
kontinuerlig	continuous,
imperium	empire,
dj	dj,
di	di,
de	the,they,
dc	d.c.,
sverigedemokraterna	sweden democrats,
stalins	stalins,stalin,
watson	watson,
människorna	men,
orolig	worried,
riktningen	direction,denomination,
du	to,you,
dr	doctor,doktor,
sattes	was added,
peyton	peyton,
offret	the victim,
runt	around,
spridningen	proliferation,the spread,
konst	art,srt,
sentida	recent,
splittrades	split,
offren	victims,
tyngre	heavy,heavier,
fågelarter	bird species,species of bird,
viktigt	important,
libanon	lebanon,
kurdiska	kurdish,
vanlig	ordinary,normal,
utförd	completed,performed,
utföra	perform,out,
förena	combine,unite,combining,
uteslutande	exclusivly,only,exclusively,
återställa	reset,resett,
präglats	been characterized,marked,
utfört	done,
massiva	solid,
utförs	out,
sexuell	sexual,
djuret	the animal,animal,
fornnordiska	old nordic,ancient nordic,old norse,
månarna	moons,
fångenskap	captivity,
piratpartiet	pirate party,
djuren	animals,
materialet	the material,material,
smaken	the flavour,flavor,
osmanska	osmanian,ottoman; osmanli,
komplikationer	complications,
we	we,
självständigheten	independence,
förkortningar	abbreviations,
miljö	environment,
jämförelse	comparative,comparison,
huvudsakligen	generally,primarily,
militären	military,the military,
garanterar	ensures,guarantees,
muhammed	muhammed,
kännetecknas	is characterized,characterized,
cox	cox,
startade	started,
kommer	is,
brad	brad,
gruppens	group (-s),
målningen	milling,the painting,
samverkan	co,cooperation,
graviditeten	the pregnancy,
kännetecken	distinction,sign,
thierry	thierry,
fångar	captures,prisoners,
chrusjtjov	khrushchev,chrusjtjov,
genomför	implement,out,
tony	tony,
slaveriet	slavery,
smith	smith,
japans	japans,japan's,
patienten	patient,the patient,
biologiska	biological,
lösning	solution,solution; resolution,
framträdande	apperance,
hitlers	hitlers,
patienter	patients,
klubblag	club team,
nära	close,
attacken	the attack,attack,
vindar	winds,
attacker	attacks,assaults,
fest	party,fest,
juridik	law,
drottningen	queen,the queen,
frekvens	frequency,
bulgariens	bulgaria,
fromstart	starting from,
vagn	carrige,
johansson	johansson,
påstådda	alleged,
kupp	kupp,coup,coup (d'etat),
aik	aik,
anhängare	supporters,
nordöstra	nordeastern,northeast,
klippa	cut,
spanjorerna	spaniards,the spaniards,spanish,
gärdestad	nugent,
have	have,
moldavien	moldova,
deltagarna	the participants,participants,
jordbruk	agricultural,
påverkades	was affected by,affected,
själva	self,actual,
våg	vague,road,wave,
patent	patent,
datorer	pc,
bergskedjor	mountain ranges,
självt	itself,
utgivna	published,
bunny	bunny,
andelen	the share,the proportion,
producerades	produced,
raid	raid,
hann	did,reached,
saddam	saddam,
balkan	the balkans,
sexualitet	sexuality,
delstater	states,
hand	hand,
delstaten	land,the state,
nervosa	nervosa,
hans	his,
bilen	the car,car,
koncentrerad	concentrated,concentration,
aspekter	aspects,
förlorade	lost,
rörelsen	movement,
kyla	cold,
riksdag	parliament; diet,the parliament,
rör	touch, move(-s),touches,
styrkorna	forces,
mamma	mother,
monaco	monaco,
rörelser	movement,movements,
röd	red,
thc	thc,
skottland	scotland,
gärningsmannen	perpetrator; offender,the offender,culprit,
newton	newton,
kall	cold,
nästan	almost,close,
kroppens	the body's,the bodies,
goda	good,
enades	agreed,
kalender	calendar,calender,
upptäckte	discovered,found,
swahili	swahili,swahilli,
lindh	lindh,
så	as,so,
distributioner	distributions,
påföljande	following,subsequent,
wright	wright,
havets	the seas,sea,
skick	state,condition,
kvinnan	woman,female,
samfund	communities,order,
plasma	plasma,
född	born,
förbättra	improve,
föda	feed,give birth; food,
återgick	returned,returning,
skadorna	injuries,damages,damage,
arab	arab,
fusion	fusion,
indianer	indians,
föds	born,
everton	everton,
engelskans	english,
hepatit	heptatitis,
acceptera	acceptable,accept,
årlig	yearly,
indelning	the subdivision,classification,
indelningen	division,subdivision,classification,
dahlén	dahlén,
xbox	xbox,
gandhi	gandhi,
transkription	transcription,transcript,
sixx	sixx,
motsvarighet	equivalent,
avsätta	unseat,depositing,
bort	away,
born	born,
presidentvalet	presidential elections,presidential election,
borg	tower,castle,
bord	table,
kungar	kings,
humor	humor,humour,
territorierna	territories,
purple	purple,
serbiens	serbias,
siffran	number,figure,
vinterkriget	the winter war,winter war,
columbus	columbus,
stadsdelarna	districts,neighborhood (-s),
vägar	roads,paths,
bevara	preserve,preserving,
fängslades	imprisoned; jailed, gaoled; incarcerated,jailed,
post	week,not a swedish word,
slovakien	slovakia,
vunnit	won,
upplösning	resolution; dissolution,resolution,
banker	banks,
ajax	ajax,
olika	different,variety,
jacques	jacques,
återfinns	found,is rediscovered,
samer	sami,
lois	lois,
epicentrum	epicentre,epicenter,
fängslade	inprisoned,imprisoned,
blivande	prospective,future,to be,
gemenskapen	the collective,community,
way	way,väg,
was	was,
war	war,
representerar	represents,
hypotes	hypothesized,hypothesis,
skiljas	separated,separate,
motorvägar	highways,
inträffar	occur,
inträffat	occurred,
partiledare	party leader,
emil	emil,
reser	travels,rise,
studierna	studies,the studies,
mtv	mtv,
finansiering	financing,
litterär	literary,
långvarig	prolonged; lengthy; long,long,
träning	training,practice,
erövra	conquer,
engagerade	dedicated,engaged,
moore	moore,
utomlands	abroad,
tesla	tesla,
xiis	xii,
efter	after,
billboard	billboard,
moln	cloudy,cloud,
empati	empathy,
toppen	the top,
cellerna	cells,the cells,
möta	meet,face,
förmåga	abilities,ability,
janukovytj	janukovytj,yanukovych,
möte	meeting,
arkitekter	architects,
test	test,
götaland	götaland,
konservatism	conservatism,
mött	met,
femton	fifteen,
tottenham	tottenham,
räknat	calculated,counted,
reglerar	regulates,controls,
regleras	is regulated,controlled,
rätter	dishes,
hemma	at home,
omgivande	surrounding,surounding,
rätten	right,the court,
solens	solar,
bergmans	bergman's,bergmans,
dance	dance,
uppfanns	was invented,invented,
tenderar	tend,
datum	date,
redaktör	editor,
osäker	unsure,
lider	suffering,suffers,
utkämpades	fought,
förhistorisk	forhistorisk,prehistorian,
afrikaner	africans,
heller	neither; nor,nor,
rådet	council,
igelkott	hedgehog,
zone	zone,
vattenånga	steam,water vapour,
terror	terror,
vänder	turn,face,
division	division,
charles	charles,
hannah	hannah,
uttrycka	express,
enskild	single,
lättare	light,easier,
hannar	males,
uttryckt	expressed,
avbröts	interrupted,
enskilt	individually,single,
salvador	salvador,
stycken	pieces; parts,pieces,
gud	god,
nedsatt	impaired,reduced,decreased; diminished,
datorspel	video game,computer game,
hisingen	hisingen,
levnadsstandard	living standard,standard of living,
frigörs	released,is released,
ljuset	the light,light,
säte	sate,seat,
formella	formal,
litterära	literary,literal,
templet	temple,
revolution	revolution,
alfa	alpha,
cosa	cosa,
engagerad	dedicated,engaged,
invandrade	immigrated,immigrant,
sköttes	operated,handled,
mål	case,mal,
formellt	formally,formal,
motsatte	opposed,
midsommar	midsummer,
stimulera	stimulate,stimulating,
motsatta	opposite,
yorks	yorks,
ungdomar	youths,adolescents,
tidig	early,
ingick	were included,was,
kosmiska	the cosmic,cosmic,
uniform	uniform,
fastigheter	real estates,properties,
utspelar	takes place,set,
syster	sister,
versionen	edition,the version,
gener	genes,
oerhörd	tremendous,
marxismen	marxism,
kärlek	love,
påstås	claimed,
klassificeras	classified,
genen	gene,the gene,
oerhört	tremendously,extremely,
tillträde	access,
antarktiska	antarctic,
flames	flames,
sistnämnda	later,last,
kemi	chemistry,
franklin	franklin,
ponny	pony,
fronten	front,the front,
vinnare	win,winner,
ekr	ekr,ad,
churchill	churchill,
marken	soil,
vapnet	the weapon,the weapon; escutheon; coat of arms; arms; badge,
spridit	spread,disseminated,
ukrainas	ukranian,ukraine's,ukrainian,
vapnen	weapons,the weapons,
krigare	warriors,warrior,
fbi	fbi,
kärnkraftverk	nuclear power plant,
presenterar	presents,present,
upprättade	established,prepared,
äktenskapet	marriage,
super	super,
territorier	territories,
stabilitet	stability,
live	live,
regel	rule,
territoriet	territory,
angels	angels,
överhuvudtaget	in general,
fransmännen	the french,frenchman,
parallellt	parallel,
club	club,
rivalitet	rivalry,
snabbt	fast,quickly,
enda	only,single,
målvakten	the goalkeeper,
zarathustra	zarathustra,
ämnena	subjects,the elements,
närmar	close,closing,close in,
varför	therefore,why,
norrköpings	norrköpings,
feministiska	feminist,
snabba	rapid,
löner	salaries,
ibm	ibm,
ibn	ibn,
interaktion	the interaction,interaction,
frukt	fruit,fruits,
can	can,cancer,
erbjuder	offers,
heart	heart,
några	few,a few,
december	december,
nobels	nobel's,
influensavirus	flu virus,influenza,
gentemot	towards,against,
abort	abortion,
uppstår	occur,
genomgått	experienced,passed,
ligan	league,
pojke	boy,
uppskattades	was appreciated,
betydelse	importance,significance,
kopplingar	connections,
perserna	the persians,
southern	southern,
riktlinjer	guidelines,
framgångarna	successes,
göteborgs	gothenburg,gothenburgs,
gräns	border,
ungern	hungary,hungaria,
förutsättning	provided,prerequisite,
romarna	romans,the romans,
flyttas	moved,
flyttar	move,
kurt	kurt,
kurs	course,rate,
ukrainska	ukrainian,
rekordet	record,the record,
maktens	the powers,forces,the power's,
landshövding	county governor,
ingripa	act,
ganska	fairly,quite,
ättlingar	descendants,
magnetfält	magnetic,magnetic field,
generalguvernören	governor general,general governor,
linnés	linnaeus,
fält	field,
skabb	mites,scabies,
idéerna	ideema,ideas,
levde	lived,survived,
utnämndes	was declared,appointed,
därifrån	from there,
bergskedjan	mountain range,the mountain group,
yngre	younger,
hals	throat,
varav	of which,which,
arton	18,eighteen,
halv	half,
nog	enough,
författarna	the authors,writers,
förvaras	stored,is stored,
komponenter	components,
begränsa	limit,
not	note,
nou	nou,
rakt	straight,
now	now,
dödsstraffet	capital punishment; death penalty,death penalty,
uppgörelse	settlement,agreement,
frihet	freedom,
språk	language,
främmande	foreign; alien,undesirable,foreign,
antyder	indicates,
stockholm	stocholm,stockholm,
januari	january,
drog	draw,pulled,drug,
aspergers	aspergers,
em	em,european championship,
el	el,
en	a,
flamländska	flemish,
ej	not,no,
ed	ed,
utbrett	wide,widespread,
spåra	track,trace,
strålningen	radiation,
ex	eg,
kroatiska	croatian,
et	et,
resultera	result,
fuglesang	fuglesang,
ep	ep,
premiärministern	prime minister,
er	you,your,
album	album,
teorier	theories,
återkommande	recurring,
videon	video,
hustrun	his wife,
kortare	shorter,
stallone	stallone,
punkt	item,point,
genetisk	genetic,
skära	carve,
välkänd	known,well-known,well known,
marina	marine,
betraktades	considered,regarded,
åt	to,
böhmen	bohemia,
british	british,
domen	judgment,verdict; judgement,
linné	linen,linneus,
allmänheten	public,general public,
arbetsgivare	employers,
blind	blind,bank,blank,
xi	xi,
förändrats	changed,
derivatan	derivative,the derivative,
ring	ring,
xv	xv,
bergqvist	bergqvist,
våglängder	wavelength,wave lengths,
omtvistat	contentious,disputed,
priser	rates,prizes,
desmond	desmond,
svenske	swedish,
sheen	sheen,
dessutom	moreover,furthermore; moreover, additionally; likewise,furthermore,
satsningar	ventures,investments,resources,
färre	less,
spelningar	tour,gigs,
fascisterna	fascists,
delats	divided,been awarded,
television	television,
europeisk	european,
sidorna	the pages,pages,
utbyggda	expanded,expand,
ändrades	changed,
kloster	monastery,
grundad	founded,based,
craig	craig,
premier	premiums,
statsminister	prime minister,
faktor	factor,
kairo	cairo,
grundat	founded,based,
grundar	bases,
grundas	is based,
anger	indicates,gives,
anges	is put at,specified,
befolkningstillväxt	population growth,befolkningstillvaxt,
hjälp	using,help,
hör	include,belong,hears,
form	form,
skär	will,cut,
fortsatte	continued,
fortsatta	continued,
etiopiska	ethiopian,etiopian,
bönor	beans,
hög	high,
online	online,
skäl	reasons,reason,
kategoriorter	category visited,
numera	now,nowadays,
santiago	santiago,
successivt	successively,progressively,
egentlig	actual; factual; real,actual,
bekostnad	detriment,expense,
dvärgar	dwarves,dwarfs,
glödlampor	lightbulbs,light bulbs,filament,
america	america,
på	on,in, on, at,
michelle	michelle,
lyfter	lift,lifts,lifting,
norrmän	norwegians,
nordligaste	northern,northernmost,
parlamentets	parliament,
runda	round,
orsaka	cause,
abraham	abraham,
skapats	was created,generated,
doktor	doctor,
kyrkorna	churches,the churches,
nazisternas	nazi,
marocko	morocco,marocco,
colombo	colombo,
teori	theory,
perfekt	perfect,
mannens	man,man's,
byggda	constructed,
rötter	roots,
varmblod	warmblood,
adolf	adolf,
raúl	raul,
himmel	heaven,
huskvarna	huskvarna,
epoken	epoch,the epoch,
dagbok	log,
sierra	sierra,
mörk	dark,
definierade	defined,
uppståndelse	resurrection,
mörker	dark,darkness,
riddare	knight,
samuel	samuel,
gudarnas	the gods',gods,god's,
ambitioner	ambitions,
folkomröstning	referendum,
marxistisk	marxist,
tävla	compete,
handlingar	actions,
drabbas	suffer,affected,
facupen	fa cup,fa-cup,
tvingade	forcing,
bushadministrationen	the bush administration,bush administration,
länge	long,
storstäder	metropolises,cities,
tillfällig	temporarily,
osbourne	osbourne,
övergången	transition,transformation,
sport	athletics,sport,
katastrofer	disasters,catastrophes,
depressionen	the depression,depression,
konstaterade	concluded,established,stated,
ladin	ladin,
depressioner	recessions,depression,
israels	israeli,israel's,
import	import,
kommunismens	communism,the communisms,
katastrofen	catastrophy,the catastrophy,
yta	surface,
ronja	ronja,
personlighet	character,personality,
flygande	flying,
männen	men,
utgivningen	the publication,the release,
verket	plant; indeed,board,
rike	kingdom,
verken	plants,wroks,
utgavs	was published,published,
comeback	comeback,
samtal	conersation,call,
monicas	monica's,
mona	mona,
bördiga	fertile,
placerad	disposed,
handlar	is,concerns,
kristinas	kristina's,crisis thawed,
propaganda	propaganda,
feminismen	feminism,
undersökning	study,
nils	nils,
comet	comet,
placerar	place,places,
placeras	placed,
utnyttja	use,
avskaffande	elimination,abolition,abolishment,
dömande	sentencing,judging,
regeringens	government,
lägenhet	apartment,appartment,
bomull	cotton,
riksrådet	riskradet,privy council; council of state; crown council; senate,privy council,
östtyska	east german,
överlever	survives,
handlande	action,
långfilm	feature film,feature movie,
oliver	olives,
välstånd	prosperity,
wien	vienna,
sker	is,
oden	node,oden,
knappt	barely,
socialdemokrater	social democrats,
dräkt	costume,outfit,
observera	note,observe,
utförda	formed,performed,made,
utförde	did,
elvis	elvis,
funnits	found,been,
ik	ik,
konservativa	conservative,
ytan	the area,surface,area,
uefacupen	the uefa champions league,
rapporter	reports,
prinsessan	the princess,princess,
rapporten	report,
polens	polands,pole,
ordningen	the order,order,procedure,
ändå	spirit,
ansikte	face,
tjeckien	czech republic,the czech republic,
eran	era,
tycker	thinks,
inslag	impact,elements,element,
finanskrisen	financial crisis,the financial crisis,
tänkande	thinking,
behandlade	treated,
kvarter	quarter,block,neighborhoods,
kenya	kenya,
västerländska	western,
katalanska	catalan,
helium	helium,
grundade	based,
infödda	natives,native,
slaget	the strike,type,
långt	far,long,
orsakade	caused,causing,
programvara	software,
media	media,
långa	langa,long,
talmannen	president,
homosexualitet	homosexuality,
kromosom	chromosome,
pesten	the plague,plague,
lite	little,a little,
figurer	figures,
speciella	special,
offensiven	offensive,
begär	requests,request,
skivbolaget	record label,the record company,
acdc	ac/dc,
omfattande	large,massive; extensive,
omfattar	encompass,include,
omfattas	comprise,subject,
speciellt	particularly,
omgående	immediately,immediate,
ekonomisk	economic,
tradition	tradition,
fredspris	peace prize,
skånes	scania,scania's,
erkänd	acknowledged,recognized,
erkänt	recognized,
flaggor	flags,
mynning	outfall,mouth,
forskarna	the scientists,scientists,
skandinaviska	scandinavic,scandinavian,
tydlig	clear,
botten	bottom,
samiska	sami,
eleverna	the pupils,the students,
lagerkvist	lagerkvist,
spänningar	tensions,
nazismen	nazism,
euron	the euro,euro,
malcolm	malcolm,
lade	laid,added,
ditt	your,
strävar	striving; aiming (to; for),strives,
irland	irland,ireland,
hovet	court,the court,
stund	while,
östergötland	Östergötland,east gothland,
selma	selma,
amy	amy,
lady	lady,
tobak	tobacco,
strävan	the quest,
nationella	national,
skilda	separate,
miniatyr|en	thumbnail,
skilde	varied,
varandra	each other,
nationellt	national,nationally,
t	t,
låga	cook,low,
astronomer	astronomers,
lågt	low,
präglades	was marked,imprinted,
stånd	position,
fönster	windows,window,
slår	switch,beats,
användbara	usable,
sålts	sold,
indikerar	indicates,
frigörelse	liberation,
berodde	depended,
agera	act,
bestämd	fixed,
strindberg	strindberg,
utskott	committee,organ,
strålning	radiation,
bestämt	decided,particularly,
nsdap	nsdap,
inuti	inside,
växa	growth,grow,wax,
kategoriledamöter	category members,category: members,
bestäms	determined,is decided,
kaffet	coffee,the coffee,
francis	francis,
övertygad	confident,
ideologi	ideology,
jamaicanska	jamaican,
central	central,center,
nordliga	northernly,northern,
socialistiska	socialistic,socialist,
sri	sri,
torget	square,
bidragen	contributions,
efterkrigstiden	the post-war period,post-war,
kapten	captain,
klassiker	classics,classic,
transporter	carriage,transports,
karriär	career,
your	your,
area	area,
specifikt	specifically,
stark	strong,
start	start,
anställd	employed,hired,
danska	danish,
specifika	specific,
likväl	nevertheless,still,
gånger	times,
fastställa	determine,confirm,
hawking	hawking,
guillou	guillou,
wailers	wailers,
sämsta	worst,
gången	time,
traditionerna	traditions,the traditions,
expeditionen	the expidition,expedition,
spänner	span,
minne	memory,
engelskan	english,
indelningar	divisions,
minns	remembers,remember,
miguel	miguel,
bilmärke	car make,
expeditioner	expeditions,
kostar	costs,
kungen	king,the king,
grammis	grammy,
sveriges	swedens,sweden,
godkände	approved,
styrde	steered,
knut	knut,knot,
transportera	transport,
nere	down,low,
mongoliet	mongolia,
efteråt	afterwards,
upphovsman	author,creator,
tänderna	teeh,teeth,
you	you,
köper	making,
knä	knee,knees,
drift	operation,drift,
översätts	translated,translate,
massachusetts	massachusetts,
röda	red,
bandmedlemmarna	band members,
skuggan	the shadow,
tjänare	servant,
handelsmän	merchants,
morgonen	the morning,am,
färdas	travels,
susan	susan,
olympiastadion	olympa stadium,olympic stadium,
monte	assembly,
eriksson	eriksson,
beskrivningar	descriptions,
energikälla	source,energy source,energy call,
messi	messi,
öknen	the desert,desert,
loppet	bore,
antoinette	antoinette,
griffin	griffin,
råvaror	raw,wood,raw materials,
lämpliga	suitable,
påbörjades	commenced; begun,was started,
lämpligt	suitable,
fästning	fortress,
skiljer	differs,is different; differ,
vers	verse,
jensen	jensen,
får	may be,can,
verk	work,works,
osv	etc.,
sanna	true,
heaven	heaven,
sverige	sweden,
behöver	need,
louis	louis,
mild	mild,
industrialiseringen	indutrialization,industrialization,
resan	the trip,journey,
uppfattas	are regarded,
rasism	racism,
magdalena	magdalena,
skiva	record,disc,
fåglarnas	the birds',birds,
egendom	property,
kritiserats	criticized,
orgasm	orgasm,
markerade	selected,marked,
trupper	troops,
utåt	outwardly,out,
stöder	supporting,supports,
tvskådespelare	tv actor,
besöker	visit,
bedrev	conducted,managed,
fjärde	fourth,
förbjuden	smoking,
erhöll	obtained,recieved,
bernhard	bernhard,
förbjuder	prohibiting,forbids,
misstänkta	suspected,suspect,
inblandad	mixed,
förbjudet	prohibited,
irak	iraq,
ersatt	replaced,
avbryta	cancel,
genomförde	carried out,
ersättare	alternate,
kronor	kronor,crowns,
observeras	observed,is noticed,
uttalat	pronounced,outspoken,
lämna	leave,supply,
uttalas	pronounced,be pronounced,
arena	arena,
medarbetare	employees,coworker,
signifikant	significant,
vår	spring,
krigen	wars,
dyker	dives,shows,
marissa	marissa,
minst	at least,
boxning	boxing,boxing; pugilism,
sagor	fairytales,tales,
kriget	the war,war,
hoppades	hoped,
perspektiv	perspective,
medicin	medicine,
då	then,when,
globen	lobe,
nazityskland	nazi germany,
gick	passed,
grunda	found,base,
dalarna	valleys,
kritiserat	criticized,criticised,
nukleotider	nucleotides,nucleotide,
familj	family,
avsedd	adapted,intended,
simba	pool,
arrangemang	arrangement,
taket	the roof,ceiling,
tillät	distillate,
etablerad	established,
förlängningen	elongation,
planen	the plan,plan,
bära	carry,mean,
oecd	oecd,
bolagets	company's,the corporation's,
representeras	represented,
expansionen	expansion,the expansion,
teatrar	theaters,
massan	mass,
kurdistan	kurdistan,
avled	died,
okänt	unknown,
utökat	extended,expanded,
blodtryck	blood pressure,
ständiga	permanent,
latinamerikanska	latin american,
site	site,
inspelad	recorded,
räknar	counts,
räknas	calculated,are counted,
lagstiftande	legislative,legislating,
ständigt	always,constant,
mördad	murdered,murderd,
företeelser	phenomena,
gazaremsan	gaza strip,the gaza strip,
ombord	onboard,board,
livslängd	life,life expectancy,
istället	instead,
trummisen	the drummer,drummer,
rapporterade	reported,
kejsardömet	empire,
partner	partner,
herrens	lord,
species	species,
ökar	increases,
gälla	valid,be valid,
serber	serbs,
ledger	ledger,
linköping	linköping,
smitta	infection,
mängden	amount,
reidars	reidars,reidar's,
ytterligare	additional,
samarbetet	co,
utför	perform,out,
long	longitude,
turkarna	turks,the turks,
torde	should,
fastän	although,
försök	experiments,expirements,
fd	former,ex,
ff	ff,
invasion	invasions,
samarbeten	cooperations,collaborations,
fn	un,the un,fn,
stabil	stable,
vattenkraft	hydroelectric power,hydro,
kostnaden	cost,
byggandet	construction,the building,
skivan	record,disc,
enzymer	enzymes,
allmänna	general,
korset	cross,
kognitiv	cognitive,
segrar	victories,
sänder	broadcast,transmits,
kostnader	cost,expenses,costs,
dream	dream,
nämnts	mentioned,above,
tillgångar	assets,
helt	completely,totally,
bloggar	blogs,
tornet	tower,the tower,
tornen	towers,the tower,
hela	entire,full,
maffian	mafia,
hell	hell,
kombinerade	combined,
eros	eros,
hundratusentals	hundreds of thousands,
romance	romance,
kompositörer	composers,compositors,
antagits	adoption,
systems	systems,system,
österrikes	austria's,austrias,
mahatma	mahatma,
musikalisk	musical,
bytte	swapped,
arsenal	arsenal,
konstitutionella	constitutional,
greps	was arrested,arrested,
dyrt	a high price,dearly,
petter	petter,
närmare	further,
fullt	full; fully; completely,completely,
fulla	full,complete,
skrivit	written,wrote,
die	die,
kontinentens	the continents,continent,
ifk	ifk,
etnisk	ethnic,
neil	neil,
positionen	position,the position,
märktes	labeled,
positioner	positions,
rättvisa	justice,
försäljning	sales,sale,
aktörer	players,actors,
robert	robert,
bodde	lived,
lungorna	lungs,the lungs,
stödet	support,the support,
pythagoras	pythagoras,
känna	known,know,
utredningen	investigation,the investigation,
heroin	heroin,heroine,
känns	feels,felt,
delningen	division,pitch,
vasas	vasa,vasas,vasa's,
svarade	answered,said,accounted (for); answered,
åtskilliga	several,
etnicitet	ethnicity,ethnic,
skogen	woods,forest,
skilja	seperate,differ; differentiate,separate,
american	american,
förbättrade	improved,
underhåll	support,entertainment,allowance,
kung	king,
skiljs	separated,separate,
sändes	was sent,sent,
utvecklats	developed,
synen	sight,
etiska	ehtical,codes,
elden	fire,the fire,
riksföreståndare	regent,
minoritetsspråk	minority language,
fabriker	factories,
helsingborgs	helsing borg,helsingborg's,
taggar	tags,thorn, twig,
synes	seems to,apparently,appears,
miss	miss,
rygg	back,dorsal,
deltagare	contestant,participants,
kanada	canada,
kongresspartiet	congress party,indian national congress,
station	station,
parlamentsvalet	parliament election,parliamentary elections,
nigeria	nigeria,
brittiska	british,
luminositet	luminosity,
brittiske	british,
delades	divided,split,
lupus	lupus,
läst	read,load,
brittiskt	british,
tvungen	forced,had,
bildande	forming,formation,
växterna	plants,
stora	large,big,
långsamt	slowly,
aristokratin	aristocracy,
andersson	andersson,
värden	values,
värdet	the value,
stiftelsen	foundation,
gren	crotch,branch,
sekunder	second,
charlotte	charlotte,
bestämdes	was determined,
teslas	teslas,tesla's,
genomgripande	radical,good,comprehensive; radical,
medeltemperaturen	median temperature,the average temperature,
tvärtom	on the contrary,contrary to,vice versa,
nominerad	nominate,nominated,
militär	military,
karl	karl,
vädret	weather,
grundarna	founders,
liberalismen	the liberalism,liberalism,
lik	similar,alike,
liv	life,
mänskliga	human,
herre	lord,master; lord,
avseenden	regard,
jämföras	comparable,compared,
mexiko	mexico,
åkte	went,relegated,
logotyp	logo,
sektor	sector,
säsongens	season,the seasons,
kan	can be,
freddie	freddie,
kap	chapter,cape,
fågel	bird,
utgör	constitutes,
himlakroppar	celestial bodies,
södra	southern,south,
förnuftet	reason,the common sense,
polacker	polish,poles,
klädd	clothed,coated,
räknade	counted,
recensioner	reviews,
rådde	prevailed,was,
två	two,
osäkra	doubtful,
ingenting	nothing,
jupiters	jupiter's,jupiter,
möjligen	possibly,
counterstrike	counterstrike,
hänvisar	reference,
muslimsk	muslim,muslim; muslem,
integritet	integrity,
justice	justice,
humanistiska	humane,humanistic,
åländska	Åland swedish,aland,
ikon	icon,
lennon	lennon,
darwin	darwin,
ingå	be a part,include,be included in,
dominans	dominant,dominance,
arabvärlden	arab world,
tillhört	belonged to,
utrikes	foreign,
gått	gone,passed,
alexander	alexander,
dogs	dogs,
restauranger	restaurants,restaurant,
avsaknaden	absence,
dömdes	sentenced,was convicted,
vilket	which,
målare	grinders,painter,
tolkiens	tolkien,tolkien's,
västkusten	the west coast,
grunden	base,
allmänt	generally,generally; public,
maurice	maurice,
bakgrund	bakground,background,
tidigare	earlier,before,
ändamål	object,purpose,
grunder	bases,
mörkare	darkey,darker,
förekom	was,
flyter	float,
direktör	director,
haddock	haddock,
pictures	pictures,
lösa	solve,
pjäser	checkers,plays,
löst	solved,dissolved,1st sentence: loosely; 2nd & 3rd: solved,
produkten	product,
chansen	chances,chance,
kategorin	category,the category,
allvar	earnest,serious,
likhet	similar,resemblance,like,
utsträckning	extent,
köket	cuisine,the kitchen,
genre	genre,
länk	link,
produkter	products,
league	league,
rankning	ranking,rating,
lejonet	the lion,lion,
anor	ancestry,lineage; ancestry,
viljan	will,te will,
slavar	slaves,
kyrkliga	religious,from the church,church,
bott	lived,
läsaren	the reader,
evolutionsteorin	theory of evolution,
uppfylla	satisfy,fulfill,
betydde	meant,ment,
derivata	derivative,
scientologikyrkan	the church of scientology,church of scientology,
linux	linux,
utgjordes	was,comprised; consisted,
sokrates	socrates,
nacional	nacional,
skydd	protection,
händerna	hands,
merparten	most,larger part,
minskade	minimum period,was reduced,
enheten	unit,
enheter	units,
oändligt	infinity,infinitely,
konsensus	consensus,
gestalt	figure,
walter	walter,
isolerade	isolated,
handlingen	the story,
budgeten	budget,the budget,
anthony	anthony,
livet	the life,life,
genomfört	carried out,carried through,
genomförs	implemented, carried through,conducted,is carried out,
socialism	socialism,
match	game,match,
hegel	hegel,
analytisk	analytical,
läser	read,are reading,
diktator	dictator,
guide	guide,
slutar	ends,end,
slutat	ended,left,
uttryckte	expressed,
nationalitet	nationality,
klippiga	rocky,
sorter	kinds,varieties,types,
bärande	wearing,leading,fundamental; wearing; supportive,
lagar	laws,
tillfällen	occasion,oppertunities,
kombineras	combined,
staffan	staffan,
kombinerat	combined,
grant	word,
borgerliga	bourgeois,conservative,
deltagande	participation,
demokratin	the democracy,democracy,
kombinerad	combined,
grand	grand,
ingår	is,penetrations,
luxemburg	luxembourg,luxemburg,
folkslag	kind of people,peoples,
kungahuset	royal family,royal house,
bon	nests,
anklagats	accused,
 km	kilometers,
kommunicera	communicate,communicating,
förlag	publishers,magazine,
seglade	sailed,
armenien	armenian,armenia,
svealand	svealand,
fatta	make,to make,
kurdisk	kurdish,
stjärnorna	the stars,
präglas	characterized,
cruz	cruz,
frihetliga	libertarian,
flygplan	aircraft,airplane,
nutid	present,
präglad	marked,characterized,
följande	following,the following,
feminister	feminists,
departement	department,
njurarna	the kidneys,kidney,
tortyr	torture,
skal	shell,skin,
fredliga	peaceful,
romerskkatolska	roman catholic,
uppfinnare	inventor,
kallblod	cold blooded,draught horse,
taiwan	taiwan,
henne	she,her,
gänget	the group,the gang,gang,
nikki	nikki,
barack	barack,barracks,
välkända	known,
varuhus	department store,
egenskap	trait,
djup	deep,
marco	marco,
bestå	consists,exist,comprise,
lika	similar,alike,
gör	does,makes,
kulturen	culture,
enklare	simpler,
kulturer	cultures,
gitarristen	the guitarist,
baserade	based,
dialekt	dialect,
läs	read,
immigranter	immigrants,
innan	before,
uppvärmningen	the warm-up,
känslig	susceptible,
releasedatum	release date,
dylikt	such,
koden	the code,code,
infektion	infection,
criss	criss,
gandhis	gandhi's,gandhi,
terminologi	terminology,
unge	young,kid,
donna	donna,
begärde	called,demanded,
tolkats	interpretation,interpreted,
kommenterade	commented,
byggnader	buildings,
biträdande	assistant,assisting,
pierre	pierre,
våldet	the violence,violence,
economic	economic,
publiceringen	the publication,publishing,publication,
syndrom	syndrome,syndrom,
sammanhängande	context of,connective,continous,
skapat	created,
världsarvslista	world heritage list,
vilda	wild,
skapar	creates,
skapas	creates,
faktorn	factor,
slash	slash,
skapad	created,
enormt	gigantic,fusionenormously,
bägge	both,
nationalistiska	nationalistic,
sarajevo	sarajevo,
run	run,
steg	rose,step,
rum	room,
sten	stone,
mellankrigstiden	interwar years,interwar period,
naturvetenskapliga	science,scientific,
offside	offside,
skrivet	written,
benfica	benfica,
bistånd	aid,assistance,
führer	fuhrer,
myndighet	authoroty,authority,
övergick	transended,went over,
linjen	line,
etablerade	established,
fysiologiska	physiological,
efterträdare	successor,
refererar	reference,
linjer	routes,lines,
edvard	edvard,edward,
länderna	states,the countries,
ändringar	changes,
ida	ida,
fåtal	a few,
stanna	stop,
egenskaper	characteristics,
ön	island,
öl	beer,
reaktorer	reactors,
semifinalen	semi finals,semifinal,
institut	institute,institution,
emellan	inbetween; between,between,
överst	top,at the top; uppermost,
föreningen	association,compound,
fokuserade	concentrated,focused,
ligga	lies, lie,lie,be,
spänningen	exitement,voltage,
består	beasts,exists,
visat	found,shown,
heritage	heritage,
spridd	spread,
jonsson	jonsson,
orsaker	causes,
ledamot	member,representative,
strukturen	the structure,structure,
japanerna	japanese,the japanese,
spektrumet	spectrum,
larry	larry,
strukturer	structures,structure,
drabbats	afflicted,
skådespelaren	actor,
skull	sake,
ute	absent,out,
nyval	re-election,election,
skuld	liability,
malin	maleic,malin,
trafikerade	frequent,trafficked,
  km²	square kilometre,km2,
politik	politics,policies,
förbjöds	banned,forbidden,
chelsea	chelsea,
ligacupen	league cup,
bränslen	fuel,fuels,
ihåg	remember,
avsåg	meant,
uppfyller	fulfills,
hårdrock	hard rock,
igenom	through,
krigets	the war's,war,
sjunde	seventh,
musikens	music,
berättat	told,
relationerna	the relationships,relations,
berättar	tells,
berättas	is told,told,
korn	korn,barley,
rester	remains,
dras	draw,preferred,
drar	drag,earn,
inkomstkälla	income cold,source of income,was added to cold,
william	william,
drag	trait; characteristic; feature,move,characteristic,
mästare	master,champion,
matematiska	mathematical,
resten	the rest,rest,
jagar	hunting,
kors	cross,
närmaste	nearest,closest,
samarbetade	collaborated,
enade	united,
medför	entails,means,
officerare	officers,officer,
tunga	tongue,
heath	heath,
tillfälliga	temporary,
folkliga	popular,folk,
tungt	heavy,
svt	svt,
dvs	d.v.s.,i.e.,
skyskrapor	high rise buildings; sky scrapers,skyscrapers,
stones	stones,
bonniers	bonnier's,bonniers,
höst	autumn,fall,
placera	position,place,
indiska	indian,
katt	cat,
företeelse	experience; phenomenon; feature,feature,phenomenon,
lutning	closing,incline,
ge	to give,give,
tänker	thinking,
ga	ga,
go	go,
gm	by,
träd	into,tree,
kate	kate,
världsrekord	world record,
baron	baron,
tillhör	belongs,belonging to,
toppar	tops,peak,
dröjde	not until,
tänkandet	thinking,the way of thinking,
wave	wave,
rinner	running,flow,flows,
kommunismen	communism,
försvarsminister	minister of defence,
michael	michael,
ryan	ryan,
utbredning	distribution,distrubution,
tidszoner	time zones,
jönköping	jönköping,jonkoping,
stift	pin,diocese,
akut	acute,
oklart	clear,
socialdemokratiska	socialists,social democratic,
zh	zh,
derivator	derivatives,derivative,
mussolinis	mussolini's,mussolini,
honan	the female,female,
geologiska	geological,
visserligen	certainly,although,
början	top,beginning,
intervjuer	interviews,
singapores	singapores,singapore's,
börjat	started,begun,
kolonialism	colonialism,
geologiskt	geologically,
mussolini	mussolini,mossolini,
kinas	kinase,chinas,
erövringar	conquests,
hansson	hansson,
bjöd	offered,invited,
polen	poland,pole,
byttes	was exchanged,
genombrott	breakthrough,
cell	cell,
experiment	experiment,
förhistoria	prehistory,
valen	elections,
gasen	gas,
utrikespolitiken	foreign policy,the foreign policy,
invigdes	inaugurated,
bindande	binding,
offentlig	public,published,
innerstaden	inner city,
händelsen	the occurence,event,
gåva	gift,
eminem	eminem,
vreeswijk	vreeswijk,
uppgick	was,
ryska	russian,
händelser	handelsar,events,
innebandy	floorball,
svenskans	the swedish language,swedish language,
västerut	west,westwards,westward; west,
chans	chances,chance,chanse,
överlevnad	survival,
förening	union,compound,
dopamin	dopamine,
uppfinningar	inventions,
avsedda	aimed,for,intended,
vuxen	adult,
italienska	italian,
genetiska	genetic,
personen	person,the person,
utdöda	extinct,
genetiskt	genetically,genetic,
kunde	could,
stärka	enhance,strengthen; bolster,
personer	person,people,
oktober	october,
sjunger	singing,
starten	start,
nordkorea	north korea,north koreans,
invigningen	inauguration,the opening,
huxley	huxley,
misslyckades	failed,
turkiets	turkey's,turkeys,
debutalbum	debut album,
släppts	released,
mottagaren	the recipient,receiver,
guds	god,god's,
kenny	kenny,
utomstående	outside people; outsiders,outside,
linköpings	linkopingas,linköpings,
halloween	halloween,
beslöt	resolved,decided,
studioalbum	studio album,
talat	spoken,spoke,
fördelningen	distribution,
talas	spoken,is spoken,
talar	speaks,speak,
romantikens	romanticism,
tåget	train,the train,
kretsar	circles,circuitry,
tågen	train,the trains,
sovjetunionen	the soviet union,
fälttåg	campaign,
ferdinand	ferdinand,
folkmängd	population size,population,
kronprinsen	crown prince,the crown prince,
oroligheter	unrest,
fara	danger,
uttalet	the pronounciation,pronunciation,
svenskar	swedish,swedes,
dödlig	lethal,mortal,
sena	late,
fars	father,
utfördes	was carried out,preformed,
ringde	called,
österrikiska	austrian,
säljer	sells,
reagerar	react,reacts,
tillhöra	belonging to,
absint	absinthe,
artisterna	artists,
encyclopedia	encyclopedia,
rörde	had something to do with,touched,was about,
kungliga	royal,
socken	parish,
högtider	holiday,feasts,
timmar	hours,
presidenter	president,presidents,
offentliga	public,
förstördes	destroyed,was destroyed,
någonting	nothing,anything,
presidenten	president,the president,
offentligt	public,publicly,
verklighet	true,reality,
belopp	amount,sum,
tränger	cut in,penetration,
begick	commited,
kyrkor	churches,
insekter	insects,
allting	everything,
filosofiska	philosophical,
naturgas	natural gas,
konserten	the concert,concert,
zagreb	capital of croatia,zagreb,
ägna	baiting,spend,devote,
läror	teachings,
front	front,
konserter	concerts,
dikt	poem,
intäkterna	the revenues,
miniatyr|px|den	miniature,
hunden	the dog,dog,
kläder	clades,clothes,
university	university,
räckte	enough,handed,
finnas	found,(be) found,
mode	fashion,mode,
förmågor	capacities,abilities,
modo	modo,
täcker	attacks,covers,
vilken	which,
föreslogs	suggested,was suggested,
usama	osama,
illuminati	illuminati,
globe	globe,
skolgång	school attendance,schooling,
 procent	percent,per,
stiger	rises,rising,
osmanerna	ottoman turks,ottomans,
apartheid	apartheid,
skov	relapse,
skor	shoe,shoes,
sandy	sandy,
endast	only,merely,
entertainment	entertainment,
förutom	besides; in addition to; aside from,except,
islamisk	islamic,
samarbetar	cooperates,collaborates,
samarbetat	collaborated,
max	max,
solsystem	solar system,
vinter	winter,
omfatta	cover,
torres	torres,
frånträde	withdrawal,
bilder	images,pictures,
lycka	happiness,good luck,
lida	sheath,suffer,
bilden	image,the image,
förstod	understood,
förbund	union,federal,league; alliance; union; compact; covenant,
kommunala	local,municipal,
livsmedel	food,
banor	paths,line,
times	times,
åter	again,undertake,
benämnas	named,entitled,
strida	conflict,fight,
tillgången	access,
tigrar	tigers,
austin	austin,
partierna	portions,
riksdagsvalet	parliamentary election,parliamentary elections,
ursprungsbefolkningen	the native population,indigenous people,indigenous population,
minoritet	minority,
brandenburg	brandenburg,
centrum	center,
bedöma	judge; decide,assessment,
kategorihedersdoktorer	category of honorary degrees,
spaniens	spain's,
ipredlagen	ipred act,
attack	attack,
boken	paper,the book,
mao	mao,
dygnet	day,
infaller	no cells,falls,
final	final,finite, final,
viktor	viktor,
belgiska	belgian,
hasch	hashish,
emellertid	however,
styrelseskick	form of government,government,
lista	list,
definierat	defined,
ben	bone,
definieras	is defined,defines,
definierar	defining,defines,
arbetade	worked,
inbördes	relative,intermutual,
israelisk	israeli,
ber	asks,
bet	bit,
julian	julian,
kvinnans	female,
hjärna	brain,
need	need,
bordet	the table,
varade	duration,
förra	last,
tredjedelar	thirds,
visor	songs,
förlorades	lost,was lost,
släkt	family,
attackerna	attacks,attack,
runorna	the runes,runes,
röst	voice,
förblev	remained,
jorge	jorge,
regn	rain,
montana	montana,
kvarstår	remains,
regi	direction,
tyskar	germans,
sändas	broadcast,be transmitted,sent,
nå	access,reach,
överföring	transfer,
skogar	forests,
långtgående	far-reaching,
platon	platon,platonic,
parker	parker,parks,
minska	reducing,reduce,
tolkien	tolkien,
fynden	finds; findings,findings,
allvarliga	severe,
försvara	defend,defending,
skedde	was,
poesi	poetry,
parken	park,the park,
hade	was,had,
basen	became,base,
baser	bases,
gemensam	common,
härskare	ruler,
förbli	remain,
varit	has been,been,
partnern	the partner,
aspekt	aspect,
psykologin	the psyhology,psychology,
boris	boris,
klassiska	classic,
inbördeskrig	civil war,
omloppsbana	orbit,
michigan	michigan,
förbjöd	forbade,forbid,
området	the area,area,
inflytelserika	influential,
klassiskt	classical,classic,
häst	horse,equine,
områden	area,
städerna	urban,
karriären	career,the career,
älskade	loved,loved; beloved,
gray	gray,
evolution	evolution,
processer	processes,
tillgång	access,
mohammed	mohammed,
grav	tomb,grave,
gran	spruce,
influensa	influenza,flu,
också	also,
grad	rate,
kvadratkilometer	square kilometers,
processen	process,the process,
vänt	turned,
sydafrika	south africa,
lätta	light,lighten,
västindien	caribbean,west india,
förband	units; formations; bound (themselves),bond,
neutralt	neutral,
korea	koreans,korea,
stats	state's,state,
tenn	tin,
individens	individual's,the individual's,
flicka	girl,
gotiska	gothic,
staty	statue,
state	state,
företagets	the company's,
ken	ken,bank,
högra	right,
ersätta	replacing,replace,
sovjetiska	soviet,sovjet,
satsa	bet,
benämningen	the designation,the name,label,
merry	merry,
jobba	work,
befälet	the command,command,
problem	problems,
hits	hits,
kaffe	coffee,
synvinkel	angle,
vulkaner	volcanos,volcanoes,
källkod	source code,
framgångsrika	successful,
trädde	met,entered,come into effect,
varierade	varied,
älskar	loves,
stratton	stratton,
framgångsrikt	successful,
partiklar	particles,
jersey	jersey,
uppsättning	equipment,set,
fördelar	advantages,share,advantage,
helsingfors	helsingfors,helsinki,
torn	tower,
opposition	opposition,
dominerande	dominating,dominant,
kategoribrittiska	category: british,category uk,
knst	knst,
leipzig	leipzig,liepzig,
johans	johan,
revolutionen	the revolution,revolution,
johann	johann,john,
kings	kings,king's,
sammanhang	connection,context,
christer	christer,
willy	willy,
trycket	pressure,
sara	sara,
fokusera	focus,
äldre	old,older,
poet	poet,
påminde	reminded,
poes	poe,poe's,
kingston	kingston,
vinci	vinci,
övertalade	over spoke,persuaded,
affärer	business,
spanska	spanish,
spanien	spain,
humör	temper,mood,
strömningar	sentiments,
kanarieöarna	canary islands,the canary islands,
 meter	meters,meter,
erbjuda	offer,
reaktionerna	reactions,
könsorganen	sex organs,the genitals,the reproductive organs,
utgjorde	made up,was,comprised; consisted of,
platons	plato,platos,
reaktion	reaction,
vilkas	whose,
rysslands	russia's,
enkel	simple,plain,
feber	fever,
demo	demo,removed,
rättigheter	rights,
mysterium	mystery,
nordirland	north ireland,northern,
måleri	painting,
kategorikrigsåret	category war years,
alfabetisk	alphabetical,
revir	turf,territory,
inre	inner,
reformationen	reformation,
parti	party,batch,
instabil	unstable,
campus	campus,
varmed	whereby,
begav	went (to),traveled,
griffon	griffon,
dickens	dicken's,dickens,
korrekta	correct,
växjö	växjö,
flygbolag	airline,carriers,
anka	anka,duck,
nationens	nation,
rankas	ranks,
särskild	specific,particular,
införa	introducing,introduce,
eklund	eklund,
nämligen	namely,
spred	spread,
alperna	alps,the alps,
lagring	storage,
flickan	the girl,
strömmen	current,the stream,
grenar	branches,
i	in,
kärleken	love,
theodor	theodor,
lugna	calm,
europarådet	european council,
onda	evil,
rösta	vote,
störta	rush,interfere,
sänds	sends,sent,
sofia	sofia,
omkom	died; was killed,died,
himmler	himmler,
förekommer	occurs,preferred is,
sända	transmitting,
sände	sent,
vida	broad,wide,
jeff	jeff,
reducera	reduce,
natt	night,
nato	nato,
sweet	söt,
titta	see,
jesper	jesper,
katolska	catholic,
utan	without,
sanning	true,truth,
vanligare	more common,
historia	history,
definitivt	permanent,
historik	history,
klassificering	classification,
loss	unstuck,off,
lincoln	lincoln,
norges	norway's,
fernando	fernando,
martin	martin,
page	page,
regeringar	rings,governments,
lager	layer,
kolonierna	colonies,
vardagliga	everyday,
pojkarna	boys,the boys,
library	library,
förlusterna	loss,
vardagligt	everyday,
förenklat	simplified,made easier,
omöjligt	impossible,
skorpan	crust,
peter	peter,
lagen	the law,law,
moskva	moscow,
skrifter	writings,
 km²	kilometres,
kaspiska	caspian,
hyser	accomodates,holds,
folkets	the people's,people,
slott	castle,
alliansen	the alliance,alliance,
fanns	was,
förde	out,
skriften	no.,writings,
broar	bridges,
hinder	obstacle,barrier,
motsättningar	oppositions,frictions; clashes,
meddelade	informed; announced,announced,stated,
samlades	collected,gathered,were united,
journal	journal,jurnal,
reza	reza,
kromosomer	chromosomes,
halvön	peninsula,the peninsula,
småland	småland,
usas	usa:s,u.s.,
keramik	ceramics,
freedom	freedom,frihet,
beslutade	resolved,decided,
samlats	collected,gathered; collected,
skrev	said,
polisens	police,
troligen	probably,likely,
synsätt	viewpoint,
hävdade	argued,claimed,
mytologi	mythology,
betydelsefulla	significant,
glenn	glenn,
underjordiska	underground,
räddade	saved,
tendenser	tendencies,
längsta	longest,maximum,
utility	utility,
hammarby	hammarby,
pc	pc,personal computer,
museum	museum,
djävulen	devil,the devil,
realiteten	de facto,reality,
afrika	africa,
distinkt	distinctive,
cricket	cricket,
north	north,
delstaterna	states,
instiftade	instituted,
neutral	neutral,
ho	ho,
behov	necessary,
hc	h.c.,
ha	be,
he	he,
samtida	contemporary,
svarta	black,
stål	steel,
fysik	physics,
allierad	ally,
dator	computer,
pippin	pippin,
komiker	comic,comedian,
förslaget	proposition,the suggestion,
hästar	horses,
invandring	immigration,
bitar	bit,pieces,
farlig	dangerous,
pelle	pellet,
ordbok	dictionary,
ibland	sometimes,
erik	erik,
själ	shawl,soul,
motsvarar	comparable,
eric	eric,
diego	diego,
omväxlande	varied,
sänktes	reduced,
närma	approach,approximate,
speciell	specific,
mineraler	minerals,
serveras	served,is served,
vulkaniska	vulcanic,volcanic,
canada	canada,
stat	state,
hittade	found,
pontus	pontus,
revolutionära	revolutionary,
musikvideor	music videos,
stad	city,
musikvideon	music video,
resulterade	resulted,
stan	town,
bly	led,lead,
hjärnan	brain,the brain,
stam	strain,tribe,
spontant	spontaneous,
etiken	ethics,
förekomma	occur,
inser	recognize,realizes,
klass	grade; class,class,
alkohol	alcohol,
blogg	blog,
konsumtion	consumption,
hinner	have time to,time,
felaktig	incorrect,error,
auktoritära	authoritarian,
protest	protest,
andra	second,
fredrik	fredrik,
flest	most,the most,
buddy	buddy,
likaså	also,as well,
upplagan	edition,
swan	swan,
kommersiellt	commercial,
kulturell	cultural,
bli	be,become,
kommersiella	commercial,
köpmän	traders,merchants,
gjordes	made,was,was made,
hemmet	the home,
kristendom	christianity,
östersjön	baltic,balticsea,
vasa	vasa,
åstadkomma	provide,create,
upplysningen	the enlightenment,enlightenment,
kända	known,
kände	felt,
examen	exam,degree,
disneys	disneys,disney,
behövdes	required,
försöka	try,
chokladen	the chocolate,
avståndet	distance,the distance,
sydväst	southwest,
nederländerna	the netherlands,netherlands,
sexton	sixteen,
dagens	current,todays,
upp	up,
rollfigurer	roll model,
force	force,
berlins	berlin,
förstaplatsen	first place,
bröstet	chest; breast,breast,
dennes	his,
avfall	waste,
neo	neo,
nej	no,
kommissionen	commission,the commission,
unescos	unesco,
ned	down,bottom,
trodde	thought,
uppdelningen	partitioning; sectionalization; division; split (-ting),splitting,division,
new	new,
representanthuset	house of representatives,
ner	bottom,
romani	romani,romany,roma,
med	with,
genomföra	perform,out,
men	but,
drev	pursued,drove,
vinden	the wind,wind,
pedro	pedro,
mer	more,
läses	read,is read,
luther	luther,
geografiskt	geographically,
därpå	then,thereon,darpa,
oro	anxiety,
åka	go,
fyllde	filled,
dubbla	double,
sju	seven,
kolonier	colonies,
geografiska	geographical,spatial,
dra	pulling,pull; (with)draw,
snabbast	fastest,
magnusson	magnusson,
reste	travelled,stood,
högtid	festival,festival; holiday,
£m	million pounds,
efterföljare	following,successors,
rosenberg	rosenberg,
reagan	reagan,
inleddes	started,began,initiated,
fördelning	distribution,
soldat	soldier,
moral	morality,
berättelserna	the stories,stories,tales; stories,
prokaryoter	prokaryote,
datorn	pc,
gävle	gävle,
lennart	lennart,
provisoriska	provisional,
bytet	the exchange,change,
oscar	oscar,
ljus	light,
nervsystemet	nervous system,the nervous system,
berlin	berlin,
upplevde	experienced,felt,
wikipedias	wikipedia,wikipedias,
ljud	noise,
köln	köln,
kategorikvinnor	category women,
flora	flora,
trots	although,
procent	percent,per,
kapitalistiska	capitalistic,
sundsvall	sundsvall,
kanadas	canada's,
erövringen	conquest,
tidskriften	the magazine,magazine,
abstrakta	abstract,
världskrigets	the world war's,world war,
förväntade	expected,
talets	the speechs,century,
klitoris	clitoris,
konstitutionen	constitution,
tusen	thousands,
tidskrifter	magazines,periodicals,
risk	risk,
sats	kit,
satt	saat,sat,
nobelstiftelsen	nobel foundation,
bonaparte	bonaparte,
avrättningen	execution,the execution,
trött	tired,
turnera	tour,
polis	police,
autonoma	autonomic,
stilla	still,stationary,
tycktes	seemed,
orsakar	causes,
orsakas	caused,causes,
orsakat	caused,
utomeuropeiska	overseas,non-european,
gård	farm,house,
könsorgan	was organ,sex organ,
klarar	do,
president	president,
orsakad	caused,induced,
indelat	divided,split,
medföra	bring,lead; result in, imply; entail,result,
indelas	divided,
indelad	divided,
medfört	resulted,led to,
låtskrivare	songwriter,
indisk	indian,
ändra	change,
kvicksilver	mercury,witty zeal,
förfäder	ancestors,
fifa	fifa,
föreställningen	the concept,show,
panthera	panthera,
ibrahimović	ibrahimovic,
munnen	the mouth,mouth,
murray	murray,
föreställningar	performances,
helena	helena,
buddhister	budhists,buddhists,
listor	lists,
personal	personal,employed,staff,
förödande	devastating,
amerikanen	american,
amerikaner	american,americans,
irans	iran's,
federationen	federation,
förstnämnda	first named,aforementioned,
aborter	abortions,
infektioner	infections,infection,
startar	begins,start,starts,
startat	started,
medlemmar	members,
downs	down,
stimulerar	stimulating,
omgivning	surroundings,ambient,
isen	the ice,
myntades	coined,was coined,
huvudrollen	the main role,leading part,
inledde	started,launched,
tillvaron	existence,life,
sida	page,side,
överraskande	surprisingly,
skeppet	the ship,nave,
side	side,
kammaren	chamber,the chamber,
bond	bond,
liga	compatible,league,
päls	fur,
mediet	medium,
medier	media,medias,
milan	milan,
aids	aids,
håret	hair,the hair,
kiev	kiev,
uppsala	uppsala,
årsåldern	age group,years old,
hänvisa	reference,refer,
talet	rate,
ihop	up,together,
talen	rate,years,
sluta	end,stop,
återfanns	was rediscovered,found,
venezuela	venezuela,
bestod	was,
foto	photo,
neutroner	neutrons,neutron,
larssons	larsson's,
normer	standards,
stöds	is supported,
nietzsche	nietzsche,
nomineringar	nominations,
uppförande	code,behavior,
folkvalda	elected,
faktum	fact,
iso	iso,
reinfeldt	reinfeld,
representant	representative,
sökte	searched,
starta	start,launch,
stewart	stewart,
gå	go,
nätet	net,
jordanien	jordan,
arrangeras	arranged,arrange,
skalvet	quake,
leddes	passed,was led,
massiv	massive,
objektet	object,
föreslagit	suggested,proposed,
girls	girls,
vikingatiden	the viking age,vikings,
förbi	past,past the,
objekten	items,the objects,
hollywood	hollywood,
någonstans	somewhere,nowhere,
representerade	represented,represent,
alfred	alfred,
åskådare	spectators,audience; viewer,
medeltiden	middle ages,
besegrades	defeated,
skaffade	acquired,aquired,
sabbath	sabbath,
grönwall	gronwall,
symptom	symptoms,
hundar	dogs,
chef	head,
formell	formal,
kontrast	contrast,
antarktis	antarctica,antarctic,
street	street,
regissören	director,
härkomst	origin,
parter	party,sides,
troligtvis	probably,
bobo	bobo,
palace	palace,
stadsdelen	the district,district,
låta	let,
mina	my,mine,
modern	modern,
självständiga	independent,sjalvstandiga,
självständigt	independent,independently,
triangel	triangle,
tecken	sign,signs,
lämnar	leaves,
lämnas	left,
lämnat	left,
der	german word,
skildringar	descriptions,
tidiga	early,
monetära	monetary,
muskler	muscles,
italiens	italy's,
tidigt	early,
tål	is resistant to,
blue	blue,
dessa	these,
bildar	serves as,form,
bildas	formed; made up (of),formed,
tåg	rail,trains,
bildat	formed,
dödsfall	deaths,
luthers	luthers,luther's,luther,
verksamma	active,
marie	marie,
typ	type,
diskuterats	been discussed,discussed,
maria	maria,
don	don,
utrustning	equipment,gear,
materiella	material,
talanger	talents,
dog	died,
slipknot	slipknot,
läsare	readers,reader,
points	point,
innersta	innermost,inner,
dos	dosage,
dop	baptism,
kristen	christian,
långvariga	long,long-standing,
koppla	coupling,connect,
införde	introduced,
hjälper	helps,shows,
västeuropa	western europe,west europe,
befälhavare	commander,
liza	liza,
droger	drugs,
skyldig	responsible,guilty,
långvarigt	prolonged,long-standing,
nevada	nevada,
odling	cultivation,
krönika	chronicle,
anländer	arrives,
folke	folke,
helhet	whole,
monica	monica,
stycke	piece,piece; part; section,
meningar	sentences,
kollapsade	collapsed,
stop	stop,
stor	big; great,large,
stol	chair,seat,
strategiska	strategic,
präster	priests,
christopher	christopher,
stod	stood,
mönster	marks,
earl	earl,
bar	bar,
bas	base,
existerar	exists,
skrivas	printed,
inlett	started,
existerat	existed,
anlades	was built,
bad	bath,
fokus	focus,
förändra	change; alter; replace,change,
gärningar	deeds,
anknytning	tie,
avvikande	different,deviant; divergent; different,
zonen	the zone,
zoner	zones,
gunnar	gunnar,
vända	turn,habituated,
dittills	thus far,so far,
vände	reversed,turned,
turnén	turn,tour,
öppnade	opened,opening,
inledningsvis	in the beginning,by way of introduction,
försvaret	the defense,repository,
naturligtvis	course,naturally,
skrift	no.,
underart	subspecies,
sorts	variety,
göta	göta,
omkringliggande	surrounding,
smguld	swedish championship gold,sm gold,gold medal in the swedish championships,
artikel	article,
armeniska	armenian,
nationalister	nationalists,
bidragande	contributors,
kämpa	fight,
motto	motto,
regelbundet	regularly,regularily,
isotoper	isotopes,
fns	un's,tris,
regering	the government,government,
näringslivet	business,industrial life,
fördraget	the treaty,treaty,
fördragen	treaties,the compacts,
kol	charcoal,coal; charcoal,
ung	young,
ernst	ernst,
regelbunden	regular,
upptäcker	discovers,discoveries,
atombomberna	atom bombs,the nuclear bombs,
mellanrum	space,gap,
nationalförsamlingen	national assembly,
synsättet	approach,view,
avsikt	intends,
interna	internal,
omstritt	controversial,
varmt	hot,warm,
basis	basis,
studerat	studied,
blodkroppar	blood cells,
cyrus	cyrus,
ting	matters,things,
frisk	healthy,fresh,
tillämpa	administer,implement,applying,
idol	idol,
centralasien	central asia,
betydelsefull	meningful,
igång	start,start up,
provinsen	province,
utseende	appearance,
sällskapshundar	pet dogs,companion dog,
namnen	names,name,
mindre	smaller,less,
etniskt	ethnic,
azerbajdzjan	azerbaijani,
blåvitt	blåvitt,bluewhite,blue and white,
etniska	ethnic,
pornografi	pornography,
paradiset	the paradise,paradise,
ix	4,the ninth,
förgäves	in vain,
albaner	albanians,
mexico	mexico,
kvinnor	female,women,
ip	ip,
sushi	sushi,
it	it,
hämnd	revenge,
cant	cant,
huvudort	main town,principal town,
im	im,
il	il,
in	in,
colosseum	colosseum,
utgåva	edition,
stoppa	stop,
konkurrensen	the competition,competitive,
vänstern	western,
framtida	future,
make	make,husband,
producerats	produced,
bella	bella,
västberlin	west berlin,
kommunistpartiets	communist party,the communist partys,the communist party,
roland	roland,
därmed	thus,therefore,
industriell	industrial,
makt	power,
benämningar	terms,names,
anglosaxiska	anglo-saxon,
atmosfären	atmosphere,the atmosphere,
försvarets	forsvarets,
övriga	others,
kim	kim,
nicklas	niclas,nicklas,
folkrikaste	populous,most populus,
akademiska	academic,
protesterna	protests,the protests,
roms	romes,roms,
vetenskaplig	scientific,
sydamerika	south america,
glädje	joy,
dåvarande	then,formerly,
värmland	wermlandia,värmland,
roma	roma,
viktiga	important,
grannländer	neighbors,neighboring countries,neighboring lander,
facto	facto,
just	right,just,
diameter	diameter,
jämför	compare,
sporting	sporting,
universitet	university,
psykos	phychosis,psychosis,
bollen	the ball,ball,
västeuropeiska	western european,
zon	zone,
human	human,
anders	anders,
beskriver	describes,
premiärminister	prime minister,
fysiker	physicist,
hävdar	states,assert,
bokstäver	letters,
troligt	likely,
hävdat	argued,claimed,
självstyrande	self-governing,independent,self-governance,
strax	soon,just,
royal	royal,
julen	julien,christmas,
memoarer	memoirs,
jules	jules,
friedrich	friedrich,
amerikas	america,
harald	harald,
borgen	castle,bail,the castle,
komintern	comintern,
språkets	the language's,language,
arkitekturen	the architecture,
gustav	gustav,
behövde	did,
kammare	chamber,
rättegång	steering wheel gang,
särdrag	feature,features,
följaktligen	consequently,
tittar	looking; viewing; viewer,
författningen	constitution,
bekräftar	confirmed,
gustaf	gustaf,
trafikeras	served,trafficked,
trafikerar	traffic,frequent,
bekräftat	confirmed,
världsdel	continent,
sjöfarten	shipping,
medborgarskap	citizenship,
kommunerna	kommunera,the municipalities,
släkting	relative,
intensiv	intensity,
litauen	lithuania,
syrien	syria,
kemiska	chemical,
vattnet	the water,
kontinent	continent,
kunna	to,be able,
dead	dead,
befolkningen	the population,population,
uppmärksammades	attention,drew attention,
jupiter	jupiter,
befann	found,located,
kemiskt	chemically,
dominerade	dominated,
tappar	drop,
statistik	statistics,
oralsex	oral sex,
kommuner	municipalities,local,
hudfärg	color,
miljöproblem	environmental problem,environmental problems,
teoretiska	theoretical,
arthur	arthur,
däggdjuren	mammals,the mammals,
säsongerna	seasons,
shakespeare	shakespeare,
hertig	duke,
filmatiserats	cinematized,been filmed,
benämns	designated,is mentioned,
knep	tricks,
angrepp	attack,
burj	burj,
versioner	versions,
bolt	bolt,
härstamma	stem,
burr	burr,
förkortas	abbreviated,reduced,
förkortat	shortened,abbreviated,
irländska	irish,
flyttat	moved,
fördelen	advantage,the advantage,
ljungström	ljungstrom,ljungström,
därutöver	addition,moreover,
maskiner	equipment,machines,
omröstning	vote,
mycket	very,much,
tillverkar	makes,
tillverkas	manufacture,
magazine	magazine,
ishockey	ice hockey,hockey,
strömmar	streams,flow,
grenen	the branch,branch,
förknippade	associated,
äktenskap	marriage,
psykisk	psychic,mental,
romantiska	romantic,
français	francais,
grundades	founded,was founded,
jens	jens,
romulus	romulus,
orsak	reason,factor,
utbildning	education,
amsterdam	amsterdam,
havsnivån	sea level,
fastlandet	mainland,
estniska	estonian,
märks	notice,labeled,noted,
tennis	tennis,
könen	the sexes,
bönder	farmers,
bolivia	bolivia,
märke	label,
hyllade	acclaimed,
själv	alone,own,himself,
norrlands	lapland's,
batman	batman,
ford	ford,
berg	mountain(-s),mountain,
japansk	japansk,japanese,
bero	depend,due,
bättre	better,
byggde	was,built,
fort	fast,quickly,
tempel	temple,
spelade	played,
positiv	positive,
slaviska	slav,slavic,
flickvän	girlfriend,
åriga	-year,
regeringen	the government,
båten	vessel,the boat,boat,
skelett	skeleton,
månens	the moon's,the moons,moon,
beteckningen	designation.........,designation,
avsnitt	section,part,episode,
phil	phil,
försörjde	living,
uttryckligen	specifically,
handelspartner	trading partner,
tosh	tosh,
kanske	may,
primtal	prime number,
byggnaden	building,the building,
vista	vista,
handen	hand,
handel	commercial,trade,
kunnat	could have been,
svärd	sword,
betala	pay,
digital	digital,
betalt	charge,
marxism	marxism,
kungamakten	monarchy,the monarchy,
ansluter	connects,
sades	said,was said,
överenskommelse	deal,arrangement,
frodo	frodo,
exporten	exports,the export,
katekes	catechism,
accepterade	accepted,
engagemang	commitment,
riktad	directed,
ökande	increasing,rising,
fss	fss,
expandera	expand,
riktat	directed,pointed,
riktas	directed (at),direct,target,
riktar	targets,target,
milt	mild,
armar	arms,
bomben	bomb,the bomb,
telefon	telephone,
spår	track,pairs,
manager	manager,
bomber	bombs,
vikingarna	the vikings,
stulna	stolen,
dä	the elder,
imperiet	the empire,empire,
avbrott	break,breaks,
uppdelning	division,partitioning,
petersburg	petersburg,
dö	die,
lissabonfördraget	treaty of lisbon,lisbon treaty,
me	me,
illa	bad,
din	yours,your,
fackföreningar	unions,
dig	up,
trenden	trend,the trend,
afrikansk	african,
anna	anna,
dit	there,where,
spets	edge; top,tip,point,
bulgarien	bulgaria,
olympia	olympia,
ville	did,wanted,
malmö	malmö,malmo,
diskografi	discography,
villa	house,villa,
slagit	held,
reklamen	the commercial,commercial; ad; advertisment,advertising,
invandringen	immigration,
rymden	space,
utlösning	release,ejaculation,trigger,
hästen	the horse,
bakom	behind,
afghanistan	afghanistan,
viktig	major,important,
kokain	cocaine,cocain,
föredrog	preferred,
bibliotek	library,
lönneberga	lönneberga,lonneberga,
somalia	somalia,
international	international,
madagaskar	madagascar,
avsluta	exit,
nationalismen	nationalism,
tibet	tibet,
henry	henry,
högkvarter	headquarters,head quarter,
avsaknad	absence,
kommun	local,municipality,
beskrivits	described,
boy	boy,
diagnoser	diagnoses,
canadian	canadian,
bor	lives,
gyllene	golden,golden; gilded,
folkmun	popular lore; popularly,colloquially,
bok	book,
mängder	amount,
extrem	extreme,
mänsklighetens	humanity's,humanities,
bolivianska	bolivian,
diagnosen	diagnosis,the diagnose,
hotell	hotel,
sporter	sports,
enorma	enormous,
utövar	carrying,exercise,
utövas	is practised,exerted,exercised,
världshälsoorganisationen	world health organization,
asiatiska	asiatic,asian,
sporten	the sport,port,
religionsfrihet	religion,religious freedom,
östasien	east asia,
platån	sycamore,the plateau,
skräck	horror,fear,
franco	franco,
hemmaarena	home ground,
tennisspelare	tennis player,
socialister	socialists,
maya	maya,
peru	peru,
kristian	kristian,
black	black,
left|px	left px,
österrikeungern	oster kingdom hungary,austria-hungary,
detaljer	details,
avsattes	deposited,dismissed,
brukade	used to,
ögon	eye (-s),eyes,
kemisk	chemical,
fartyget	ship; vessel,boat,
fly	escape,
hända	may,
hände	happened,
tokyo	tokyo,
mästarna	the champions,
söka	search,searching,
träffades	met,was met,reached; met,
vittnen	witnesses,
akademien	the academy,academy,
präglade	characterized,
anslutna	connected,
bristande	wanting,lack,
sökt	pending,
ulf	ulf,
hiroshima	hiroshima,
crazy	crazy,
kenneth	kenneth,
uruguay	uruguay,
winston	winston,
agent	agent,
bemärkelse	meaning,sense,
skadades	was wounded,damaged,
council	council,
dennis	dennis,
kunglig	royal,
pink	pink,
diskuterades	discussed,
oslo	oslo,
engelsmännen	english people,the english,the british,
varor	products,
ekonomiska	economic,economical,
till	to,
gitarrist	guitarist,
nya	new,
nye	new,
mat	food,
regeringstid	term of government,term of government; term of office,
överensstämmer	conform,agree,
uppföljare	sequel,
fotboll	football,
läkare	doctors,doctor,
maj	may,
upphört	ceased,left the association,end,
man	is,one,
asien	asia,
johnson	johnson,
kulturella	cultural,
sådana	such,
eng	eng.,
tala	speaking,speak,
block	block,
basket	basketball,
romantiken	romance,romanticism,
undantag	exception,except,
sådant	such,
lsd	lsd,
bussar	bus,
bevisa	prove,
alfabetet	alphabet,the alphabet,
unionen	union,the union,
gällde	applied,applied to,was,
sällsynta	rare,
moralisk	moral,
huvudsak	in principal; chiefly,main thing,
lyrik	poetry,
motståndet	the resistance,the resistence,
verksam	active,effective,
landskap	province,landscape,
juryn	jury,
sekter	sects,
inkomster	income,
äkta	married,genuine,
nazisterna	nazis,
policy	policy,
växte	grew,
main	main,
texas	texas,
lägst	lowest,lowermost,
steget	step,
kräver	requires,
janeiro	janeiro,
domstolar	courts,
försörjning	sustentation,supply,
sibirien	siberia,
leds	passed,
vindkraft	wind power,
färg	colors,colour,
uppskattning	appreciation,estimated,
leda	lead,
villkoren	the terms,conditions,
rock	rock,
föremål	object,subject,
tysklands	germany's,germanys,
guevara	guevara,
latin	latin,
tacitus	tacitus,
hellre	rather,more preferably,
söner	sons,
vattendrag	water,streams,watercourse,
avkomma	progeny,offspring,
girl	girl,
dianno	di'anno,dianno,
saudiarabien	saudi arabia,
enastående	exceptional,outstanding,
jackson	jackson,
håkansson	hakansson,håkansson,
avrättningar	execution,
pamela	pamela,
områdena	the areas,
tronföljare	heir,heir apparent,successor,
kattdjur	felidae,cat,
valdes	representatives',selected,chosen; elected,
premiären	premiere,premier,
ansiktet	face,
monster	monsters,
ort	neighborhood,place,location,
konstnär	artist,
chiles	chiles,chile's,
tomt	empty,blank,
inriktade	oriented,
california	california,
miley	miley,
brooke	brooke,
kognitiva	cognitive,
ord	word,
tunnelbanan	subway; tube; underground,the subway,metro,
keith	keith,
verkade	appeared to,were active, worked, was active,
gott	good,practically; good,
anledning	reason,
preventivmedel	contraceptives,
självmord	self-killing,suicide,
uppvisar	shows,
rankningar	ranking,rankings,
vision	vision,
stängdes	closed,
kraftig	strong,
first	first,
centrala	central,
grupperna	groups,
intryck	appearance,
uttalanden	statements,
här	this; here,is,here,
rachel	rachel,
folklig	popular,folk,
lat	methacrylate,
centralt	central,centrally,
skapandet	creation,the making,
kommunism	communism,
grundämnet	the element,element,
missnöje	dissatisfaction,
homogen	homogenous,
visar	is,shows,
visas	shown,
västbanken	the west bank,westbank,
grundämnen	elements,
individ	individual,
örebro	Örebro,
öronen	lugs,the ears,
besluten	decisions,
anus	ass,anus,
köpenhamns	copenhagen,copenhagen's,
fysiska	natural,physical,
fysiskt	physically,physical,
danny	danny,
löstes	solved,dissolved,
drevs	concentrated,was driven,
beslutet	the decision,
konkreta	specific,
fiender	enemies,
fienden	enemy,the enemy,
medlemmarna	members,the members,
lugn	calm,
jordytan	earth's surface,earth crust,
fordon	vehicle/-s,vehicles,vehicle,
inträde	entry,
marklund	marklund,
jämlikhet	equality,
stadsdelar	districts,city districts,neighborhoods,
marijuana	marijuana,
större	greater,bigger,
formerna	forms,
tänder	teeth,
orsakerna	the causes,
kevin	kevin,
adeln	nobility,
nikola	nikola,
politiska	politic,political,
förälskad	in love,
menas	mean,
skulptur	sculpture,
centralbanken	centralbank,central bank,
potential	potential,
politiskt	political,
performance	performance,uppträdande,
centralstation	central station,
magnetiska	magnetic,
channel	channel,
riktningar	direction,direction (-s),
norman	norman,
normal	normal,
morden	murders,
dagbladet	dagbladet,
halvan	half,
politisk	political,
teoretiskt	theoretic,theoretical,
mordet	the murder,murder,
arbetat	worked,
civilisationer	civilizations,
visades	was,
otaliga	countless; endless,countless,
lojalitet	loyalty,
drottning	queen,
grammatik	grammar,
österut	eastwards,
kontrolleras	is controlled,controlled,
kontrollerar	controls,controls; controlling,
ungdom	youth,
civilisationen	civilization,
show	show,
adolfs	adolf's,adolf,
regioner	regions,
or	or,
generalsekreterare	the secretary-general,secretary general,
samlingsalbum	compilations,
helig	holy,
dick	dick,
historier	stories,history,
passande	fitting,suitable,matching,
historien	history,
statsmakten	the government,power,government,
karolinska	caroline,
experimenterade	experimented,
ges	given,be given,
ger	gives; is giving,give,gives,
raser	races,
klasser	classes,
kulturellt	culture,cultural,culturally,
konsolen	bracket,
motsvarande	corresponding to,corresponding,
skådespelare	actor,
inspelningarna	recordings,
personliga	personal,
vintergatan	milky way,the milky way,
firade	celebrated,
ledaren	leader,conductor,
gen	gene,
beskyddare	protector,patron,
himmlers	himmlers,himmler,
mattis	mattis,
bengtsson	bengtsson,
statistiska	statistical,
tsaren	the czar,czar,
spridda	spread,scattered,
europacupen	euro (-pean) cup,european cup,
london	london,
tolfte	twelth,twelfth,
relativt	relative,relatively,
sämre	poor,
sekulära	secular,
fokuserar	focuses,focus,
toppade	topped,
relativa	relative,
sean	seab,sean,
slöt	closed,
utgiven	published,
menat	meant,
menar	mean,means,
kandidater	candidates,
försvarsmakten	national defense,armed forces,
döden	death,
vanns	was won,
människan	man,people,
söndagen	sunday,
personligt	personal,private,
erövrades	conquered,concoured,
människas	human's; man's,human,
landets	the country's,its,
förenta	united,
august	august,
ju	the,
tur	turn,tour,
forskaren	researcher,
jr	jr.,junior,
åker	go,treats,field; going,
timme	hour,
tum	inch,inches,
fick	got,was,
signaler	signals,
lexikon	lexicon,
kirsten	kirsten,kristen,
ministrar	ministers,
rugby	american fotboll,rugby,
ån	on,from,the river,
utvalda	selected,selected; chosen,
tour	tour,
paret	pair,the couple,parathyroid,
ås	ridge,
år	the year,year,
vätska	fluid,liquid,
tryck	press,print,
vilja	will,like,
århundraden	centuries,
cancer	cancer,
statschefen	the head of state,head of state,
syntes	synthesis,
grundare	founder,
territorium	state,
mätningar	measurements,measurments,
ryggen	the back,back,
barry	barry,
överföra	transmit,transfer,
bildats	formed,
ja	yes,
industrin	industry,
västliga	western,
utsatta	exposed,
mars	march,
överförs	is transferred,
plötsligt	suddenly,
marx	marx,
mary	mary,
kultur	culture,
flaggan	flag,
cobain	cobain,
partido	partido,
avskaffa	abolish,
bmi	bmi,
dvärghundar	miniature dogs,
spelfilmer	motion pictures,feature film,feature films,
klädsel	cover,
meningen	sense,
fortsatt	further,continued,
sound	sound,
metall	metal,
dragit	dragged,preferred,
uppstod	developed,was,
kategorimän	category: men,category men,
insåg	realized,
nionde	ninth,
sahara	sahara,
intressanta	interesting,of interest,
uppmanade	urged,encouraged,
liknande	similiar,similar,
sydkorea	south koreans,south korea,
hålls	maintained,maintaned,is held,
par	pair,
upplagor	editions,
jesu	jesu,
edwin	edwin,
same	lapp,
hålla	hold,keep,
röka	smoking,
stött	met,supported,
pan	pan,
samt	also,as well as,
tidvis	times,
hösten	fall,the fall,the autumn,
running	running,
kuba	cubans,cuba,
teknisk	technical,
lösningar	solutions,
sömn	sleep,
fattas	taken,
bang	bang,
wahlgren	wahlgren,
identifiera	identification,
gates	gates,
münchen	munchen,munich,
bebyggelse	settlement,settlements,
privatliv	private,
reaktionen	reaction,
dinosaurierna	dinosaurs,dinasaurs,
skapelse	creation,
väst	west,the west,
byggnad	building,
reaktioner	reactions,
våld	violence,force,
jakten	the hunt,hunt,
ideologiskt	ideologically,ideological,
grannländerna	neighbors,
bowie	bowie,
livstid	lifetime,life span,
programledare	host,
gotland	gotland,
ideologiska	ideological,
motverka	counteract,
trä	wood,
möter	meets,
vintern	the winter,winter,
schwarzenegger	schwarzenegger,
underarten	subspecies,sub species,
mån	concerned,
mor	mother,
haft	had,
prägel	character,mark,
mot	against,
kategori	category,
jakt	hunt,hunting,
temperatur	temperature,
mon	mon,
underarter	sub-species,subspecies,
baltiska	baltic,
kollektiv	collective,public,
mod	courage,mod,
christina	christina,
adams	adams,
födda	born,
började	started,began,
födde	gave birth too,born,
jordbävningar	earthquakes,
manhattan	manhattan,
mänsklig	human,
sågs	observed,was observed,
göran	göran,request,
bipolära	bipolar,
göras	be made,be made through,
rikskansler	chancellor,
kategorisveriges	category sweden,
feodala	feudal,
maos	maos,mao's,
förs	out,led,rapids,
jordbruket	the agriculture,
lotta	raffle,
fört	lead,
sudan	sudan,
reportrar	reporters,
föra	pre,
före	ahead (of), before,present,
ända	as far as,up,
demokratisk	democratic,
traditionell	traditional,conventional,
samman	together,
moderata	moderate,moderates,
vistas	present,
tunnlar	tunnels,
londons	london's,
framstående	prominent,
olof	olof,
akon	akon,
tongivande	influential,
tillverka	producing,
sjätte	sixth,
celler	cells,
island	iceland,icelandic,
allians	alliance,
metaforer	metaphores,metaphors,
lands	land,on land,
lagarna	the laws,
retoriken	rhetoric,
herbert	herbert,
kort	short,
arvid	arvid,
wilde	wilde,
beskrivas	described,be described,
einstein	einstein,
mark	ground, soil, territory,ground,
intellektuella	intellectuals,intellectual,
floderna	floods,rivers,
fullständigt	full,
gravid	pregnant,
behandling	treatment,
varelse	creature,
emellanåt	once in a while,occasionally,
anfalla	attack,
välmående	healthy,well-being; affluent,prosperous,
fullständiga	full,complete,
kvinnlig	females,female,
tillfälligt	temporarly,temporary,
eget	own,
inletts	started,initiation,
utbredd	widespread,spread,
birger	birger,
härifrån	from here,here,
e	e,
egen	own,
woman	woman,
tävlingen	competition,contest,
vhs	vhs,
exemplar	copies,example,
bibliografi	bibliography,
manuel	manual,
verkliga	real,fair,
identifierade	identified,
humanismen	humanism,
parlament	parliament,
håkan	håkan,
följde	followed,
youtube	youtube,
manliga	male,
öns	the islands,island's,
prestigefyllda	prestigious,
skriven	written,
palats	palace,
arabiska	arabic,arabian,
goebbels	goebbels,geobbels,
film	film,
diktaturen	dictatorship,
again	again,
genrer	genres,
effekt	effect,power,
istanbul	istanbul,
spåren	the tracks,wake,
rubiks	rubiks,rubik's,
muren	wall,
produktiv	productive,productivity,
stannade	stayed,
spåret	groove,
genren	genre,
faktorer	factors,
däremot	on the contrary,however, on the contrary,however,
ordna	arranging,arrange,
profet	prophet,
ungarna	the kids,kids,the young,
förändrade	changed,
rykten	rumors,
ledning	conduit,guidance,
henriks	henry,
kyros	cyrus,
världsliga	worldly,
kväll	evening,
nöjd	content,
palestinska	palestinian,
uppfostran	upbringing,
medicinskt	medical,
kuwait	kuwait,
snabbaste	rapid,fastest,
begå	commit,
resolution	resolution,
åtskilda	separated,separate,
mellanöstern	middle,the middle east,
vila	rest,
socialismen	the socialism,socialism,
dollar	dollar,
vill	will,to,
hindrar	prevent,stop; prevent,prevents,
ingripande	negative,intervention,
inspirerad	inspired,
liam	liam,
levern	the liver,liver,
sund	healthy,sane,
symbolen	the symbol,
kategorilevande	category of live,
rwanda	rwanda,
symboler	symbols,
skydda	protection,
skriver	write,type,
seriens	series,
kasta	discard,throw,
avhandling	treatise,thesis,
handlade	was (about); traded,was,
israeliska	isrealic,
fall	where,
ramen	frame,
stödja	support,
kulminerade	culminated,
miljoner	millions,
båtar	boats,
bröderna	brothers,the brothers,
suttit	been,sat,
ockuperades	occupied,
cornelis	cornelis,
massor	lots,tons,
växthuseffekten	the greenhouse effect,
intressant	interestingly,of interest,
material	material,materials,
abc	abc,
danmark	denmark,
abu	abu,
östtysklands	osttysklands,
public	public,
lärare	teacher,
värderingar	evaluations,values,
långhårig	rough,long haired,
bebott	inhabited,
närhet	close,closeness,
vald	selected,
jonas	jonas,
free	free,
benen	legs,
valt	chosen,selected,
sångare	singer,
historiker	historians,
jackie	jackie,
airport	airport,
uppslagsverk	encyclopedia,
alexandria	alexandria,
sjukhuset	hospital,
africa	africa,
nacka	nacka,
släktingar	relatives,
varianterna	variants,the diversities,
rösterna	votes,
författaren	the author,author,
hyllning	tribute,tribute; homage,
eye	eye,
medlem	member,
torrt	dry,
utmärkelsen	award,the award,
budskapet	message,
innebar	was; meant; entailed,was,
utmärkelser	commendations,awards,
torra	dry,
landet	state,the country,
diamond	diamond,
människa	human,man,
romersk	roman,
koma	coma,
brist	non,failure; lack of,
tillkommer	reside,will be,
hundraser	breed of dogs,breeds,
skivor	plates,records,
berätta	tell,
vladimir	vladimir,
länkar	links,
des	des,
det	is,
roosevelt	roosevelt,
utsläpp	emission,emissions,
bron	bridge,the bridge,
del	part,
lindgren	lindgren,
den	it,
lagerlöf	lagerlof,
befintliga	current,existing,
samtliga	all,
hastigt	rapidly,fast,
latinets	latin,the latin,
sovjetunionens	soviet union's; soviet's,soviet union,
betoning	stress,
hjälpte	helped,
sjukdom	illness,
medförde	resulted,brought,
födseln	birth,the birth,
sträng	string,strang,
robinson	robinson,
protein	protein,
makten	power,the power,
hämta	retrieve,fetch,
stil	type,
psykotiska	psychotic,
georgien	georgia,
stig	stig,path,
verkligheten	real,reality,
sammanfaller	coinciding,coincides,
försvinner	disappears,disappear,
primära	primary,
vikten	importance,weight,
makter	powers,
hoppade	jumped,
avtalet	the contract,
pettersson	pettersson,
laboratorium	laboratory,
ännu	even,yet,
judiska	jewish,
huvudkontor	central office,headquarters,
ligger	is,
vatten	water,
rastafarianer	rastafarian,rastafarians,
rockgrupper	rock bands,
facebook	facebook,
paz	paz,
konservatismen	conservatism,
civila	civil,
inåt	inwards,inwardly,
uppgav	said,
nordsjön	north sea,
officiella	official,
latinamerika	latin america,
fältet	the field,field,
förmågan	the ability,
göra	do,do; doing,
mörkt	dark,
gradvis	gradually,progressively,
tvåa	second,
lava	lava,
mörka	dark,
görs	is,made,is made to,
officiellt	official,officially,
människans	humans,mankinds,human,
längden	lenght,
diskussion	discussion,
ärftliga	genetic,
edmund	edmund,
inbördeskriget	civil war; civil war,civil war,
andré	andre,
odlade	grew,cultured,
saknades	missing,
trossamfund	religious communities,
suverän	terrific,sovereign,
good	good,
träffar	meets,hits,
ställas	set,be set,prepared,
planerna	the plans,plans,
fängelse	prison,
sexuellt	sexual,
oxford	oxford,
skrifterna	scriptures,
association	association,
toronto	toronto,
robbie	bobbie,robbie,
kungarna	the kings,kings,
namibia	namibia,
byggt	building,built,
anslöt	joined,
trådlös	wireless,
house	house,
energy	energy,
hard	hard,
flytta	move,
byggs	building,
förenade	united,
energi	energy,
seder	subsequently,custom,
perry	perry,
sanningen	truth,the truth,
östman	Östman,
sällsynt	rare,
oftast	usually,most often,
infrastrukturen	infrastructure,
ölet	the beer,beer,
forskning	research,
perro	perro,
förföljelser	pursuits,persecutions,
fullständig	full,complete,
konflikt	conflict; strife,conflict,
prins	prince,
lawrence	lawrence,
strömning	flow,
eventuella	any,
blekinge	blekinge,
uralbergen	urals,
eventuellt	eventually,possibly,
viken	gulf,
helsingör	helsingor,elsinore,helsingör,
inflationen	inflation,
investeringar	investments,
finland	finland,
jordens	earth,
demokratiska	democratic,
utöver	addition,
fått	was given,with,
styre	governance,rule,
legenden	legend,
ensam	alone,
styra	controlling,steer,
top	top,
sjunkande	sinking; decreasing,decreasing,
dont	do,
säkerhetsråd	security,security council,
treenighetsläran	doctrine of the holy trinity,trinity,school of trinity,
snarast	rather,as soon as possible,
juridiska	legal,
carter	carter,
förklarade	explained,said,
kom	came,
diskriminering	discrimination,
gator	streets,
kon	group,
åtta	eight,
observationer	observations,
förhindrar	prevents,prevent,
kategoriasiens	category of asia,
costa	costa,
kardinal	cardinal,
järnvägar	failways,rail,
triangeln	triangle,the triangle,
part	party,
gudarna	the gods,
domstolen	court,the court,
direkta	direct,
matteusevangeliet	gospel of matthew,
följden	the cause,result,
b	b,
avtal	agreement; deal,agreement,contract,
proteinerna	proteins,
ö	o,
personens	person,the persons,
börjar	starts,starts to,start,
hellström	hellström,
baháí	baha'i,bahá'í,
avtar	declines,avatar,
självständig	independent,independently,
följder	impact,consequences,
följdes	followed,was followed,
rikedom	riches,
försökte	try,tried,
bränsle	fuel,
gjord	made,
flertalet	most,majority; plurality,
gjort	made,done,
mountain	mountain,
hundratals	hundreds of,hundreds,
svagare	weaker,weak,
infrastruktur	infrastructure,
caesar	caesar,
genast	at once,immediately,
taktik	tactic,strategy,
inkomsterna	revenue,
dramatiskt	dramatic,dramatically,
skjuta	delay,postpone; shoot,
militärt	military,
patterson	patterson,
krafter	forces,
gillade	liked,approved; liked,
niclas	niclas,
kraften	the force,
utbrott	outbreak,outbreaks,
samtidigt	while,
organiserade	organized,
högt	high,highly,
ko	co,cow,
km	km,kilometers,
kl	at,
kr	kronas,
liechtenstein	liechtenstein,
organisk	organic,
organism	organism,
thomas	thomas,
venedig	venice,venedig,
kvalitet	quality,
bergman	bergman,
relation	ratio,relation,
utveckla	developing,
fina	beautiful,fine,
nämns	mentioned,
antagit	adopted,presumed,
konto	account,sign,
kristna	christian,
undre	lower,
wallenberg	wallenberg,
medverka	take part,participate,
världens	the world,the worlds,
tionde	tenth,
religionerna	religions,
förbudet	ban,the union,
avseende	regard,for,
blomstrade	flourished,
typiskt	typically,typical,
nationalpark	national park,
beyoncé	beyoncé,
beslutar	decides,
vänskap	friendship,
express	express,
beslutat	resolved,
förklarat	explained,declare,
typiska	typical,
förklarar	explains,
gamla	ancient,old,
husen	housing,the houses,
skickas	is sent,
skickar	sends,
brukar	usually,used to,
boende	resident,accommodation,
gamle	old,
uttrycket	the expression,expression,
uttrycker	express,expressing,express (-es),
flykt	escape,
huset	housing,the house,
svarar	responds,
somrar	summers,
stadium	stage,
styrdes	governed,
suveränitet	sovereignty,
rollfigur	character,
godkännas	approved,be approved,
höglandet	the highland,
tengil	tengil,
fann	found,
rovdjur	predator,
fans	fans,
landsbygden	rural,rural area,
champagne	champagne,
romarriket	roman empire,the roman empire,
bildandet	formation,establishment,
professionella	professional,
framförs	is presented,performed,
framfört	expressed,
rörelserna	the movements,movement,
kritiserades	critisized,critizised,
framföra	express,convey,
skivorna	records,
marilyn	marilyn,
musklerna	muscles,the muscles,
statligt	state,governmental,
uppfattning	understanding,view,
praktiskt	convenient,
statliga	state,
restaurang	restaurang,restaurant,
baltimore	baltimore,
romska	romani,roma,
beta	graze,beta,
globala	global,
kroatiens	croatia's,croatias,
förklaring	explanation,statement,
point	point,
folkmord	genocide,
karaktären	character,
andas	breath,breathes,
karaktärer	characters,
således	hence,thus,
tennessee	tennessee,
globalt	globally,global,
behöll	kept,retained,
försäljningen	sales,
lyfta	lift,
våningar	floors,storeys,
laos	laos,
bestämde	determined,chose,
inför	before,
bengt	bengt,
popularitet	popularity,
gav	gave,
effektiva	effective,
gas	gas,
vana	familiar,used,
kalmar	kalmar,
effektivt	effective,
trupperna	troops,the troops,
detsamma	the same,same,
bild	picture,image,
motorväg	freeway,highway,
åtalades	was charged,was prosecuted,
spridning	diffusion,distribution,proliferation,
bill	car,
döptes	renamed; named,renamed,baptised,
portugal	portugal,
arenan	arena,the arena,
elektronik	electronics,
påbörjade	started,
monroe	monroe - it's a persons name,monroe,
rederiet	the shipping company,shipping company,
dödat	killed,
granska	examining,
sjuk	disease,
dödar	kill,kills,
dödas	killed,
hamna	end,
motståndaren	the opponent,adversary,opponent,
administrationen	administration,
dödad	killed,
tyder	indicates,
sittande	fitting,
development	development,
övertogs	were taken,overtaken,
skotska	scottish,
syd	south,
konstnärliga	artistic,
syn	sight,view,
jerusalems	jerusalem's,
moment	step,
kallades	was called,called,summoned,
parentes	brackets,
avsett	avset,intended,
nämnde	mentioned,said,
småningom	eventually,
tillbehör	accessory,
nämnda	said,
kungariket	kingdom,
noll	zero,
kapitel	chapter,
albanien	albania,
jorderosion	earth erosion,soil erosion,
ministerrådet	minister counsellor,ministers,
skott	shots,
albanska	albanian,
norrland	norrland,northern,
dikter	poems,
bibeln	bible,
kommunister	communists,
juventus	juventus,
halvt	half,
organization	organization,
verkställande	executive,
passerar	passes,pass,
struktur	structure,
senaste	last,
alternativt	alternatively,alternative,
analytiska	analytical,
alternativa	alternative,
tropisk	tropical,
sektion	section,
kubas	cuba's,cuba,
administrativt	administrative,administratively,
monarkin	monarchy,the monarchy,
dömd	sentenced,convicted,
administrativa	administration,administrative,administative,
åtal	prosecution,
bin	bin,
dubbelt	double,
bil	car,
teknik	technic,
big	big,
kejsaren	emperor,the emperor,
avlidna	diseased,deceased,
af	of,
möttes	met,
bit	piece,
indonesiska	indonesian,
planeterna	planets,the planets,
rené	rene,
grå	gray,grey,
kolonialtiden	the colonial times,colonial period,
princip	principle,principal,
möjlig	possible,
brett	broad,
stränga	severe,
kristina	kristina,
tillstånd	state,to the dental,condition,
anatomi	anatomy,
google	google,
identisk	identical,
egyptiska	egyptian,
tolkningar	interpretations,
back	reverse,
historisk	historic,historical,
studerar	study,studies,
cocacola	coca cola,coca-cola,
lars	lars,
västergötland	västergötland,
flygplatser	airports,
måste	have to,must,
lasse	lasse,
per	per,
pratar	talks,talking,
självstyre	autonomy,self-governance,self-government,
energin	the energy,energy,
lösningen	the solution,solution,
därför	because,therefore,
nordamerika	north america,
resande	travelers,travelling,
vasaloppet	vasaloppet,
påven	the pope,pope,
ockuperade	occupied,
britannica	britannica,
korta	short,
värmestrålningen	heat radiation,
uppfattningar	opinions,perceptions,
fallit	fallen,fall,
jimmy	jimmy,
grammy	grammy,
styrelse	government; direction,board,board of directors,
barcelonas	barcelona,
steven	steven,
ordnar	decorations,
brita	brita,
ontario	ontario,
framträdde	appeared,emerged,
ökningen	increase,
ansvar	responsibilities,
turkiska	turkey,turkish,
medvetande	consciousness,consciousnesses extensive,awareness,
lyssnar	listens,listen,
jaga	course,hunt,chase,
serie	comic; row; succession; serial,cartoon,series,
konsul	consul,
bostäder	residences,housing,
torsten	torsten,
jonathan	jonathan,
skillnaden	the difference,
ledningen	conduit,the lead,
mångfald	diversity,variety,
planet	planet,
smycken	jewlery,
sultanen	sultan,
planer	plans,
amfetamin	amphetamine,
skillnader	differences,
reggaen	reggae,
jordbävningen	earthquake,
reidar	reidar,
titel	title,
expedition	caretaker,expidition,expedition,
förbjudna	forbidden,prohibited,
hjärnans	brain,
tropiskt	tropical,
tropiska	tropical,tropic,
materia	matter,materia,
tyskland	germany,
västerås	vasteras,västerås,
voltaire	voltaire,
familjer	families,
årstiderna	seasons,the seasons,
familjen	the family,family,
betalar	paying,pay,
makedonien	macedonia,
anser	view,
anses	be,deemed; regarded,
konspirationsteorier	conspiracy theories,
lena	lena,
utvecklade	oral,
länders	countries',countries,
samla	collecting,collect,
mutationer	mutations,
nådde	reached,
ritualer	rituals,
storkors	the grand cross,
talades	spoken,spoke,
regionala	regional,
sambandet	the connection,connection,
dramatiker	playwright,dramatist,dramatists,
judisk	jewish,jew,
sorg	grief,
regionalt	regional,regionally,
at	at,
flod	basin,river,
uppgår	is,
jason	jason,
stänga	close,off,
stred	fought,
uran	uranium,
frankrike	france,
förut	requires,
sigmund	sigmund,
övergav	abandoned,
intensivt	intensive,hard,
privat	private,
lilla	small,
tillämpningar	applications,implementations,
landslaget	the national team,team,
betrakta	view; regard,view,
sydafrikanska	south african,african,
sahlin	sahlin,
konsten	art,the art,
intensiva	intensive,
kollaps	collapse,
atlas	atlas,
graven	the grave,grave,
passiv	passive,
luleå	luleå,
kampanjen	campaign,
plikt	duty,
släppte	released,
tjänade	earned,
varnade	warned,
färöarna	the faroe islands,
nonsporting	non sporting,
svts	svts,
tävlingar	competitions,contests,
exemplet	the example,example,
knight	knight,
joel	joel,
ände	end,
slutade	quit,ending,
madeira	madeira,
warszawa	warsaw,
naturens	nature's,nature,
joey	joey,
förlust	loss,
störtades	overthrown,
överhöghet	supremacy,suzeranity,
utbredda	widespread,spread,
vanligaste	frequent,
cellen	cell,the cell,
påsken	easter,
höjdpunkt	climax,high point,
carlo	carlo,
depression	depression,
sträcker	stretches,extend,
går	is,goes,
chicago	chicago,
spåras	trace,
tillkomst	origin,established,advent,
senare	latterly; later,later,
sauron	sauron,
placering	position,placement,
börje	börje,borje,
analsex	anal sex,
och	and,
kyrka	church,
öar	islets,islands,
extremt	extremely,extreme,
ordförande	chairman,
börja	start,
extrema	extreme,
isländska	icelandic,
befolkningstäthet	population density,the population density,
populäraste	rated,most popular,
störning	noise,
honom	his,him,
svårigheter	difficulties,
medeltid	medieval,
turkar	turks,
alaska	alaska,
lagts	added,
katolicismen	catholisism,catholicism,
lagförslag	bill,lagforslag,
miljard	billion,one billion,
klassisk	classical,classic,
honor	ära,
färgade	colored,
existens	existence,
protokoll	protocol,
uppnår	achieve,reaches,
uppnås	obtained,is achieved,
talare	speakers,spoke,
privata	private,
stundom	sometimes,somtimes,
når	reach,reaches,
nås	reached,is reached,
filippinerna	filipinos,the philippines,
betraktas	considered,
betraktar	regard,sees,
ovan	above,
lima	lima,
somrarna	the summers,summers,
skivbolag	record label,record company,
kinesisk	chinese,
skotsk	scottish,
chi	chi,
gruppspelet	group stage,group play,
fånga	capture,capturing,
nobel	nobel,
döpt	baptized,
söder	south,
nytta	good,useful,
geografisk	geographic,geographical,spatial,
titanics	titanic's,titanic,
konkurrens	competition,
prinsen	prince,the prince,
ledamöterna	commisioners,the members,
förstå	understand,understandable,first,
utropade	exclaimed,cried out,
bakterier	bacteria,
självständighet	independance,independence,
avsikten	purpose,
iii	iii,
platsen	place,site,
ansvaret	responsibility,
britney	britney,
tunnel	tunnel,
gabriel	gabriel,
påbörjas	start,starts,
halt	content,stop; level,stop,
baserad	based,
kedja	chain,
kategorisvenska	category: swedish,
baseras	based,based on,
baserar	base,based,
baserat	based,
kyrkan	the church,church,
väldet	empire,violence,the rule,
fotosyntesen	photosynthesis,
titlar	titles,
do	do,
mozarts	mozart's,mozart,
förlängning	overtime; extension; prolongation,extension,
cecilia	cecilia,
fett	fat,
democracy	democracy,
internationellt	international,internationally,
lanserade	introduced,launched,
hendrix	hendrix,
internationella	international,
tjänst	service,
vilhelm	vilhelm,
revs	described,was demolished,
böckerna	books,
rousseau	rousseau,
riktig	real,
klar	clear,done,
trycktes	was published,printed,
föddes	was born,
herrlandskamper	herrlandskamper,men's international contest,
brändes	burned,burnt,
spannmål	grain,cereals,
förbundskapten	manager,
klan	clan,
gammal	old,
terrier	terrier,
siv	siv,
finländska	finish,finnish,
rådhus	town hall,courthouse,
dryck	beverage,drinks,
förekommit	occurred,
billboardlistan	billboard list,bilboardlist,
grannar	neighbors,
registrerade	data,noted,
olyckan	incident,
alltjämt	remains,
omslaget	cover,the cover,
dy	younger,
halvklotet	hemisphere,
strid	conflict,fight,
georg	georgian,georg,
innebär	means,
industrier	industries,
le	le,
människor	human,
la	la,
variationer	variations,
berget	mount,the mountain,
föreställer	depicts,
tillägg	addition,appendix,
weber	weber,
dag	day,
spektrum	spectra,spectrum,
utfärdade	issued,
slags	kind,type,
dam	dam,lady,
dan	dan,
valet	selection,the election,
avslöjar	reveals,
tillkommit	been,accured,
periodiska	periodic,
das	das,
sammanhanget	connection,context,
installera	installing,
day	day,
kontinuerligt	continuous,continous,
beslut	decision,
morris	morris,
newtons	newton,newton's,
syftade	alluded to,aiming,
emo	emo,
lysande	brilliant,illuminating,
engelskspråkiga	english-speaking,the english language,
juridisk	legal,
krita	chalk,
humanism	humanistic,humanism,
pitts	pitts,
kristiansson	kristiansen,kristiansson,
dokumentär	documentary,
inspirerade	inspired,
segern	victory,
programmet	program,the application,
arbetskraft	workforce,labor,
fattigdomen	poverty,
nödvändiga	necessary,essential,
matt	dull,
jerusalem	jerusalem,
mats	mat's,attention,
kärnan	core,the core,
nödvändigt	neccessary,necessary,
deras	their,
försäkra	make sure,
red	eds,
återta	retake,regain,
filmatiseringen	film version,
roterande	rotating,
frank	franks,
webbplats	website,site,
franz	franz,
odlas	cultured,
arbetare	workers,
ronald	ronald,
längre	longer,
josé	jose,
fart	off,speed,
efterträddes	succeeded,
medelhavsområdet	mediterranean,the mediterranean region,the mediterranean area,
referenser	references,
farbror	uncle,
fotografier	photographs,
nivå	level,
south	south,
liberaler	liberals,
stämmer	correct,
genomgår	undergoes,undergoing,
pga	due,
uppges	reported,
uppger	states,state,
innehålla	include,contain,
insikt	recognition,
levnadsstandarden	the standard of living,living standard,standard of living,
fruktade	feared,
omständigheter	event,circumstances,
veckan	weeks,the week,
leder	leads,leading (to),
utlopp	outflow,outlet,
energikällor	energy resources,sources of energy,
kantonerna	cantons,
förklara	explain,declaring,
maidens	maidens,
leden	hinge,lines,the route,
palestina	palestine,
demonstrationer	demonstrations,
bundna	tied,bonded,
släktet	the genus,
stället	instead,the place,
ställer	running; causing,set,
innehade	held,possessed,
firades	celebrated,was celebrated,
pågående	current,ongoing,
sjögren	sjögren,
ledamöter	commissioners,
släkten	genera,the family,
ställen	spots; places,places,
bevarats	protected,preserved,
beskrivningen	description,
domaren	judge,the judge,
matematisk	mathematical,mathematic,
inne	inside,
sweden	sweden,
kvalificerade	qualifying,
universum	universe,
mälaren	mälaren,
premiär	prime,premiere,
havs	at sea,sea,
aristoteles	aristoteles,aristotle,
tids	time,
operativsystem	os,
följd	following,
älgar	moose,
följa	follow,
basist	bassist,
uganda	uganda,
idag	today,
rådande	prevalent,
följt	followed,
följs	followed,
låt	let,
mil	mile,swedish miles,mil,
min	my,
mia	mia,
fötter	feet,on its feet,
kroppar	bodies,
tidningar	press,magazines,
mig	me,
mix	mix,
låg	low,
experter	experts,
besättningen	crew,
lån	loan,
konstverk	work of art,artworks,
konkurrerande	competing,
kommunikationer	communications,
resurser	resources,
resultatet	the result,result,
dinosaurier	dinosaurs,
varandras	each others,each other,
missionärer	missioners,missionaries,
resultaten	the results,results,
sedan	then,since,
sist	finally,last,
efternamn	last name,lastname,
liknade	looked like,similar,
stranden	shore,
upprustning	renovation,
irakkriget	iraq war,
republikanska	republican,
rörelsens	movements,movement,
milano	milano,
deuterium	deuterium,
tidskrift	newspaper,magazine,
capita	capita,
definiera	defining,define,
viktigaste	most important,
styrka	strength,power,
utgångspunkt	starting point,point of departure,
obelix	obelix,
text	text,
komplicerad	complicated,
existerande	current,existing,
inhemsk	domestic,native,
ugglas	owl,ugglas,
fungerade	thought,working,
kurfursten	elector,
rumänska	romanian,
järnvägen	railroad,rail,
euroområdet	eurozone,euro area,convergence report,
rytmiska	rhythmic,
satan	satan,
shahen	the shah,shah,
säker	items,safety,
bryssel	brussels,
organiska	organic,
snitt	on average,average,
arean	the area,area,
förändrades	changed,
buddhismen	buddhism,buddism,
överlägset	far,
förstår	understand,forstar,
regimen	regime,
studenterna	students,
uppehåll	residence,pause,hiatus,
richards	richards,
från	from,
vinsten	the win,gain,
organ	body,organ,
županija	country,
nazitysklands	nazi germany's,nazi germany,
vinster	gains,
majoriteten	the majority,
lyckade	successful,
byggdes	was,was built,
ronaldo	ronaldo,
militärer	military,
krävdes	were required,
national	national,
svenska	swedish,
eleonora	eleonora,
kapitalet	capital,
svenskt	swedish,
först	first,
bön	nests,prayer,
debutalbumet	the debut-album,debut album,
reform	reform,
redan	has already,
konverterade	converted,
intog	seized,occupied,took,
carlsson	carlsson,
avslutades	closed,ended; concluded,
vänta	(have to) wait; expect,
bör	live,should,
terräng	terrain,off,
ordentligt	properly,firmly,
översikt	overview,over term,
koncept	concept,
industrialisering	industrialization,
uppskattade	estimated,appreciated,
listan	the list,
hårdare	harder,tougher,
säkerheten	the security,safety,
översättas	translated,be translated,
viktigare	important,more important,
läsning	read,
hämtade	taken,brought,
buddhas	buddha's,buddhas,
empathy	empathy,
miniatyr|karta	thumbnail map,miniature|map,
återförening	reunion,
litteratur	literature,
aktuellt	current,relevant,
kommunicerar	communicates,
kröntes	crowned,
aktuella	current,
kommendör	commandor,commander,
förekomst	presence,
sachsen	sachsen,saxony,
fester	celebrations,parties,
inneburit	meant,resulted,
befogenhet	warrant,authority,
utsågs	was,was appointed,
medicinsk	medical,
elektroner	electron,
news	news,
ad	ad,
västmakterna	western powers,
tunisien	tunisia,
grupperingar	groups,grouping,
slippa	avoid,
gaza	gaza,
igen	recognize,back,
define	define,
asteroider	astroids,asteroids,
jämna	even,
genomsnittlig	average,
stationen	station,
stationer	stations,
orange	orange,
deep	deep,
uppmärksammat	attention,noticed,
an	an,
napoleon	napoleon,
augusti	august,
bruket	use,the use,
kraftiga	strong,powerful,
stalin	stalin,
ar	is,
ocheller	and/or,
betraktade	watched,
externa	external,
kväve	nitrogen,
tagits	taken,
flyktingar	refugees,
betalade	payed,paid,
fördrag	agreement,treaty,
vistelse	stay,
prosa	prose,
utom	except,out,
händelserna	the events,events,the happenings,
lämnade	did,left,
wolfgang	wolfgang,
blodtrycket	the blood pressure,blood pressure,
sångerna	song are,the songs,
omedelbart	immediately,immediate,
heinrich	heinrich,
hinduismen	hinduism,
kallad	called,
kontrollera	control,controlling,
framförallt	above all,in particular; above all,
kallat	called,
kallas	called,
kallar	call,calls,
center	center,
öde	fate,
seth	seth,
antonio	antonio,
sett	seen,
hoppas	hope,
omgångar	in turns; periods; mandates,cycles,
svensk	swedish,
undvika	prevent,avoid,
position	position,
deltar	part,participates,
stores	great,the great's,
kontaktade	contacted,
passade	suiting,suited,fit; suited,
mystiska	mysterious,mystical,
wagner	wagner,
misshandel	assault,abuse,
grekiskans	greek,
flertal	several,majority group,
bevarade	preserved,
vanligt	usual,normal,
hamburg	hamburger,
kampf	kampf,
reformer	reformers,reforms,
anhöriga	relatives,kin,
lake	lake,
mentala	mental,
landområden	land areas,land,
streck	bar,
belgrad	belgrade,
förnuft	reason,
uppmärksamhet	attention,attantion,
uppträder	occur,performs,
dubai	dubai,
demens	dementia,
innehöll	containing,
tusentals	thousands,
viruset	virus,
likt	like,
journalist	journalist,
works	works,
uppträda	appear,occur,
gudomlig	divine,
albumets	album,album's,
starkaste	strongest,the strongest,
värmlands	varmlands,värmlands,
etablerades	established,was established,
minsta	minimum,
est	est,
joachim	joachim,
katarina	katarina,
löser	solve,
skildrar	depicts,portrays,
skildras	is depicted,depicted,
gisslan	hostages,
internationalen	international,
definitionen	the definition,
nattetid	overnight,
definitioner	definitions,
starkare	strong,stronger,
leopold	leopold,
arterna	the species,species,
about	about,
socker	sugar,
ärkebiskopen	archbishop,
glada	happy,
mäktigaste	powerful,
slutgiltiga	final,
andel	percentage,share,
anden	spirit,
folkräkningen	census,
värd	host,worth,
alexanders	alexanders,
förstärka	strengthen,enhance,
kapital	capital,
omgiven	surrounded,
potatis	potato,
monarken	the monarch,monarch,
chris	chris,
ljusare	lighter,
föredrar	prefer,preferred,
vimmerby	vimmerby,
hatar	hate,hates,
ridge	ridge,
densamma	the same,same,
skog	wood,forest,
kuben	cube,the cube,
strävhårig	hispid,wirehaired,
föga	little,hardly; little,
flyg	flight,airforce,
kärnor	core,
medicinska	medical,
klockan	clock,o'clock,
civilbefolkningen	civilian population,the civilian population,civilians,
ryssarna	russians,
brand	fire,
bröder	brothers,
ersättning	replacement,
flygvapnet	air force,
kraft	force,power,
bud	bid,bids,
araberna	arabs,
vetenskap	science,
utrymme	space,
arbetsgivaren	employer,
lissabon	lisbon,
australiens	australia,australia's,
nedre	lower,bottom,
innanför	inside,
minuter	minutes,
vänstra	left-hand,left,
hästens	horses,horse's,horse,
circus	circus,
paraguay	paraguay,
tolkningen	interpretetation,interpretation,
omloppsbanor	orbits,
autism	autism,
betydande	important,significant,
vinner	gaining,wins,win,
manlig	male,
identitet	identity,
särskilda	special,
proteinet	the protein,
proteiner	proteins,
einsteins	einstein,once a,einsteins,
uppfattar	percieves,interpret,
picchu	picchu,
stimulans	stimulation,stimulating,
betonade	emphasized,
out	out,
försämrades	decreased,worsening,
uppfatta	perceived,perceive,
sjön	lake,
tämligen	rather,fairly,tamil again,
astronomi	astronomy,
variation	diversity,variety,
koncentrationsläger	concentration,concentration camp,concentration camps; kz-camps,
akademisk	academical,academic,
ärkebiskop	archbishop,
cirkel	circular,
philips	philips,
fakta	fact,
winnerbäck	winnerback,
baker	baker,
svag	weak,
uppfattningen	comprehension,view,
framför	in front of,particularly,
förbundet	the union,association,
okänd	unknown,
nelson	nelson,
mäktiga	powerful,
brottslingar	criminals,
slogs	fought,was,
båt	boat,
resor	travels,travel,
påsk	easter,
arkitekt	architect,
antisemitiska	antisemetic,antisemitic,
ozzy	ozzy,
granskning	review,
anfallet	the attack,attack,
upphör	end,
paris	paris,
tillväxten	growth,
deltagit	part,participated,
kapacitet	capacity,
under	for,under,
läge	mode,
svårare	difficult,
nordost	the northeast,northeast,
pommern	pommern,pomerania,
ägande	owning,
jack	jack,
invånare	resident (-s),
evert	everted,evert,
ovanstående	above,
tagit	taken,
utmärks	characterized,
utmärkt	excellent; superb; marked by; characterized by,excellent,
öppna	open,
plural	plural,
venus	venus,
matematik	mathematic,mathematics,
verklig	real,
reklam	advertising,advertisement,
parten	party,
markerar	selects,
kropp	body,
bönderna	farmers,
manus	script,
läget	location,
indierna	indians,
läger	camp,
stridigheter	oppositions,strife,
aktivt	active,
drivande	drive,driving,
ebba	ebba,
notera	note,
liberty	liberty,
aktiva	active,
zink	zinc,
kub	cube,
disney	disney,
egyptens	egypt,egypts,
språken	languages,
prata	talk,
flera	multiple,
medelhavsklimat	mediterranean climate,
utredning	study,investigation,
beck	beck,pitch,
parlamentariska	parliamentary,
preparat	substance,
studio	studio,
rysk	russian,
sommartid	summer-time,summer,during summer,
komplex	complex,komplex,
studie	study,
språket	language,
forum	forum,
lagras	stored,
ty	for,
precis	precisely,exactly; precisely,just,
proportioner	proportions,
svante	svante,
gällande	current,regarding,
koloniserades	is colonized,colonized,
upptäckter	discoveries,discovery,
upptäcktes	discovered,
julie	julie,
erektion	erection,
julia	julia,
övers	transl,
nazistiska	nazi,
hittades	was found,
misslyckats	failed,
upptäckten	the discovery,discovery,
försvarsmakt	armed forces,
eftervärlden	posterity,the world,
volym	volume,
mattias	mattias,
klassas	classified,
vinst	profit,win,
miniatyr|px|en	miniature,
konserterna	the concerts,concerts,
västtyskland	west germany,
skicka	send,
behandlingar	treatments,
romaner	novels,
växt	plant,
återstående	remaining,
muse	muse,
övertala	convince,persuade,
ludvig	louis,ludvig,
ansökte	applied,
världsarv	world heritage,
fermentering	fermentation,
rörelse	movement,
belgiens	belgium,belgium's,
igelkottens	the hedgehog's,hedgehog,
henri	henri - it's a name,henri,
mm	millimeter,
arméns	the army's,arm,army's,
antiken	the ancient world,antiquity,
ms	motor ship,
mr	herr,mr,
johanssons	johansson,
avstå	desist,
utgick	started,
partiets	the party's,parties,
ghana	ghana,
sträckan	distance,the distance,
utlöste	triggered,
persien	persia,
trädgård	garden,
florida	florida,
djur	animals,
genomfördes	was,was carried out,
fröken	miss,
ena	one,
end	end,
smält	melted,
iiis	iii's,3's,
väpnade	armed,
ens	even,
gata	street,
elektriskt	electric,
elizabeth	elizabeth,
beskrev	depicted,described,
målen	cases,goals,
förståelse	understanding,
mest	most,mostly,
västvärlden	west,western world,
målet	target,the target,
miniatyr|px|ett	miniature,
elektriska	electrical,
frågade	asked,
 cm	centimeters,cm,
nagasaki	nagasaki,
kategorier	categories,
kubanska	cuban,
galilei	galilei,
beteenden	behavior,
kontrollen	control,the control,
existera	exist,
beskrivit	described,
praxis	practice,
arbetar	work,works,
kejsare	emperor,
kampen	the fight,fight,
over	over,
arresterades	was arrested,
vitt	white,widely,
besittningar	holdings,possessions,
synonymt	synonymously,
frivillig	optional,
vita	white,
expansion	expansion,
bibelns	the bibel's,the bible's,bible,
brinner	on fire,burns,
evans	evans,
edith	edith,
nytt	new,
statschef	head of state,
dött	dead,died,
blott	merely,only,
historiens	historys,
dem	those,
senast	last,
produktion	production,
upptagen	busy,occupied,
avskaffandet	elimination,abolition,abolishment,
ansvarar	charge,
alex	alex,
jämförelser	comparison,
detroit	detroit,
ersattes	was replaced by,replaced,
ställdes	prepared,
newport	newport,
storlek	size,
ursprungligen	initially,originally,
växter	plants,
önskemål	requests,demands,
gymnasium	high school,
group	group,
dessförinnan	before (that),before,
träffade	met,
innehållande	containing,
platina	platinum,
nio	nine,
medelålder	middle age,
behövs	required,is needed,
god	good,
receptorer	receptors,
användningen	use,the use,
ammoniak	ammonia,
hemland	homeland,
riktning	direction,
danmarks	denmarks,denmark's,
paulus	paulus,paul,
got	got,
behöva	need,
independence	independence,
smala	narrow,
snuset	snuff,
icke	non,none,
herman	herman,
värnplikt	military service,
kandidat	candidate,
fred	peace,
statsöverhuvud	head of state,
undervisade	taught,
samlade	collected,
inom	within,in,
drygt	good,approximately,
statsministern	prime minister,head of state,
studera	study,
tolerans	tolerance,
bredvid	beside,next to,
vetenskapliga	scientific,
samhälle	society,
befolkade	populated,
vetenskapligt	scientifically,scientific,
transporterar	carrying,transports,
transporteras	is transported,
nyheter	news,
säsong	season,
museet	the museum,museum,
museer	museums,musser,
föreslagits	suggested,was suggested,
nhl	nhl,
institutioner	institutions,
rikaste	the richest,richest,
tillåts	is allowed,allowed,
yngsta	youngest,
sexuella	sexual,
nyheten	news,
mercury	mercury,
vikingar	vikings,
tor	thu,
yngste	youngest,
punkten	point,
merkurius	mercury,
å	on,
konventioner	conventions,
ton	tonne,tone,
punkter	points,seq,
tom	tom,
uppkommit	generated,arisen,
tog	was,took,
fördes	sea were entered,out,
adjektiv	adjective,adjectives,
ifrågasatts	is questioned,questioned,
livealbum	live album,
skildes	separated,was seperated,
meddelande	message,
rädsla	fear,
fördel	advantageously,advantage,
kulturarv	cultureheritage,cultural heritage,
territoriella	territorial,
dramer	plays,
slutsats	conclusion,
mjölk	milk,
uppmuntrade	encouragement,encouraged,
bridge	bridge,
rad	range,line,
nedgång	decline,decreases,fall,
tänka	thinking,think,
rak	straight,linear,
somliga	some,
störningar	interruptions,disorder,
växer	growing,grows,
ras	race,ras,
adhd	adhd,
övervikt	obesity,
tycks	appears,
tänkt	expected,supposed; intended,
ray	ray,
industriellt	industrially,industrial,
hittats	found,
kvällen	the evening,evening,
situationer	situations,
jorden	earth,earth; earth; underground,
lanseringen	the release,launch,
användning	use,use; usage,
öarna	the islands,
industriella	industrial,
academy	academy,
situationen	situation,the situation,
mekaniska	mechanical,
grundskolan	elementary school,
tvingas	forced,system,
skepp	vessel,ship,
elektricitet	electricity,
fralagen	fralegen,the fra law,
motsatt	opposite,
framgångsrik	successful,
motsats	contrary,
tanzania	tanzania,
metal	metal,
sekt	sect,
metan	methane,
sjöar	lakes,parks,
inflytande	influence,
agnes	agnes,
utkanten	the outskirts,outskirts,
dyrare	more expensive,expensive,
idrott	sport,sports,
saga	saga,story,
järnvägarna	the railways,railways,
queen	drottning,
gränserna	borders,limits,
radio	radio,
earth	earth,
sagt	said,
radie	radius,
absolut	absolute,absolute; total,
skada	damage,
claude	claude,
florens	florence,florens,
vinna	win,
institution	institution,
ägare	owner,owners,
gods	domain,goods,
holländska	dutch,
publik	audience,public,
återstår	remains,remain,
andras	others,
länder	countries,
mängd	amount,laden,
kommunisterna	communists,communist,the communists,
guatemala	guatemala,
gogh	gogh,
haiti	haiti,
sträckor	distances,
ålder	age,
stadskärnan	town/city,
taubes	taubes,
ändras	be changed,change,
ändrar	changing,change,
ursäkt	excuse,apology,
ändrat	changed,modified,
lovat	promised,
publicerades	published,
tidningen	the newspaper,journal,paper,
utvisning	penalty,expulsion,
kroppen	body,the body,
sakta	slowly,
ockuperat	occupied,
fördomar	bias,prejudice,prejudices,
kristendomen	chritianity,christianity,
utformade	formed,
behålla	container,keep,
mur	wall,
brinnande	burning,
antikens	ancient,
populär	popular,
slottet	castle,the castle,
finger	finger,finder,
förstås	course,mean:,
allra	very,most,-most; most,
mun	mouth,oral,
herding	herding,
förhållande	in relation,ratio,
ordnade	arranged,parent,
betonar	emphasize,
omvänt	vice versa,
maniska	manic,maniac,
seden	the seed,custom,
dödsorsaken	cause of death,
bildriksdagsval	image election,
nummer	number,
store	great,
kreativitet	creativity,
autonomi	autonomy,
anfall	attack,
verka	operate,appear,
lösningsmedel	solvent,
läggs	is,put before; submitted; put,
farliga	dangerous,
allierades	allied's,allied,
begränsade	restricted,
förbränning	combustion,
avgöra	determine,decide,
lägga	put,add,
november	november,
hitler	hitler,
solljus	sun light,sunlight,
skapades	generated,created,
rumänien	romania,
reglera	expell,controlling,
möjliggjorde	made possible,allowed,
därefter	thereafter,
hastighet	speed,
diktatorn	the dictator,dictator,
homosexuell	homosexual,
skalan	scale,
öster	east,
modernare	mor modern,more modern,
anspråk	claim,
spritt	spread,
drömmar	dreams,
invasionen	invasion,the invasion,
älgen	elk; moose,moose,
n	n,
petrus	petrus,
schizofreni	schizophrenia,
depp	depp,
förståelsen	the understanding,
claes	claes,
della	della,
nationer	nations,
viking	viking,
darwins	darwin,darwins,
därigenom	by which,thus,thereby,
vojvodskap	voivodships,voivodeship,
brott	breach,crimes,
anlände	arrived,
känsliga	susceptible,1st&2nd: fragile 3rd: sensitive,bilge accordance,
nationen	the nation,
kartan	the map,map,
vanföreställningar	delusions,
varefter	whereafter,
ekonomin	the economy,economy,
ernman	ernman,
äger	owns,
pekar	pointer,pointing,
erhållit	obtained,received,
ökade	increased,
ersatte	substituting,
pekat	pointed,identified,
negativ	negative,
welsh	welsh,
hundra	hundred,one hundred,
formatet	the format,size,
ersatts	replaced,
återvände	returned,returning,
återvända	return,
uppsving	boost,
gudom	deity,
dylan	dylan,
generna	genes,the genes,
charlie	charlie,
spelad	played,
tillkännagav	announced,
svavel	sulfur,
kemikalier	chemicals,
fattigare	poorer,
louisiana	louisiana,
jean	jean,
spelat	played,
spelas	played,
spelar	gaming,
mytologin	mythology,
kraftigt	heavily,
järn	iron,kon,
ämnen	agents,
torah	torah,
graden	rate,
europaparlamentet	the european parliament,european parliament,
grader	degrees,
picasso	picasso,
utföras	be,performed,
kolväten	hydrocarbons,the hydrocarbon,
kalifornien	california,
använt	using,used,
värnpliktiga	conscripted,inductees,
gavs	was,gave,
belagt	coated,
eld	fire,
grundaren	the founder,founder,
aktiv	active,
rätta	correct,come to grips; court; correct,
regionerna	regions,
enlighet	according (to),according,
nobelpriset	the nobel prize,
benämning	term,name,title,
donau	danube,donau,
ämnet	substance,subject,
tillgänglig	available,provided,
protesterade	protested,
auktoritet	authority,
omvärlden	world,surrounding world,
gift	married,
såväl	both,as well as,
ladda	load,
modersmål	native language,
bosnienhercegovina	bosnia-hercegovina,
specifik	specific,
tillåtna	allowed,
fotbollen	soccer,
hund	dog,
gifter	marries,toxins,
lagstiftningen	law-making,legislation,
enat	united,
hanhon	he/she,male-female,
hushåll	household,
besöka	visit,
jennifer	jennifer,
malaysia	malaysia,
donald	donald,
besökt	visited,
saturnus	saturn,
skapa	create,creating,
estetik	aesthetics,
ultraviolett	ultraviolet,
totalt	total,complete,wholly,
användare	users,
gösta	gosta,
icd	icd,
diktatur	dictator,dictatorship,
utse	appoint,name,
totala	total,
karaktäriseras	characterizes,is characterised,
elitserien	elite series,elitserien,
monoteism	monotheism,
ishockeyspelare	hockey player,ice hockey player,hockey players,
tillbringar	spends,
män	males,men,
spelare	player,
hotellet	the hotel,hotel,
meyer	meyer,
titeln	the title,
tvingades	forced,had,
systrar	sisters,
omgången	round,
plus	plus,
internationell	international,
tydliga	clear,obvious,
genomslag	impact,breakthrough,
primitiva	primitive,
skrevs	written,was,
civil	civil,civilian,
menade	meant,said,
systemet	the system,system,
tydligt	clear,obvious,
isberg	ice berg,iceberg,
sinne	mind,
anorexia	anorexia,
oförmåga	inability,failure,
omges	surrounded,
omger	surrounding the,
lagt	laid,added,
kjell	kjell,
sicilien	sicily,
gia	gia,
metabolism	metabolism,
wittenberg	wittenberg,
dialekterna	dialects,
fadern	the father,
skulden	the guilt,
barrett	barett,barrett,
fängelsestraff	imprisonment,prison,
italien	italy,
skulder	debts,liabilities,debt,
finns	there is,
eventuell	any,
fusionen	merger,
säkerhet	safety; security,
amerikanerna	americans,the americans,
värvade	recruited,referred,
tillika	also,well,
araber	arabs,
behandla	treatment,
trio	trio,
bildt	bildt,
bilda	form,
läsa	read,
tronen	throne,the throne,
kambodja	cambodians,
förbud	ban,prohibiting,
liberalism	liberalism,
tätorten	conurbation,agglomeration,
ni	you,
margareta	margareta,
no	no.,
tillverkade	manufactured,made,
when	when,
nf	nf,
finna	found,
ny	new,
tio	ten,
lösas	solved,
nr	no.,number,no,
tätorter	urban,conurbation,
nu	now,
picture	picture,
phoenix	phoenix,
sätts	is,is placed,
miscellaneous	miscellaneous,
gäster	guests,
tunna	thin,
massakern	massacre,
sätta	insert,set,
kronprins	crown prince,
väckte	awakened,aroused,
beroendeframkallande	addictive,
vietnam	vietnam,
cellens	cell's,
rom	rome,rom,
ron	ron,
rob	rob,
rod	rod,
dvärg	dwarf,
roy	roy,
koreanska	korean,
udda	odd,
fiktiv	fictitious,
laura	laura,
mottagarens	the reciever,the receivers,
konstitutionell	constitutional,
bär	carryng,berries,here,
tanke	light,in light of,
federation	federation,
även	also,
läns	county,
varvid	in which,
underhållning	entertainment,
flytt	escaped,move,fled,
krossa	crush,crushing,
metod	method,
inlärning	learning,
brother	brother,
christmas	christmas,
olyckor	accidents,
lever	living,liver,
tillverkningen	production,the production,
församling	congregation,assembly,
införandet	introduction,the introduction,
trend	trend,
stilar	styles,
kategorirock	category:rock,
linda	winding,linda,
colin	colin,
svartån	svartån,
förorter	suburbs,
port	gate,port,
uppgifterna	data,
ifråga	with regards to,challenged,
passa	match,
agnosticism	agnosticism,
miniatyr	miniature,thumbnail,
ögat	eye,
cykel	bicycle,cycle,
månaderna	months,
angelina	angelina,
gräs	grass,
gravitation	gravitation,gravity,
kamp	struggle,fight,
vindkraftverk	wind turbine,
enkla	simple,single,
metaller	metals,
eiffeltornet	the eiffel tower,
jord	earth,
turister	tourists,
dublin	dublin,
sina	their,his,
införts	been inserted,introduced,
lokal	local,
ankomst	arrival,
filmen	the movie,film,
tilltagande	increasing,
rafael	rafael,
luften	air,
sikt	term,run,
etablera	establish,up,
trummor	drums,
bolaget	company,the company,
ungerska	hungarian,
russell	russell,
undan	escape,
utropades	proclaimed,was proclaimed,
samfundet	association,
lp	lp,
anda	spirit,
inblandade	involved,
andy	andy,
kurder	kurds,
australian	australian,
turné	tour,
crüe	crüe,
uppskattningar	estimates,
typerna	the types,
staten	state,
kär	in love,
övergå	transition,transend,
palestinsk	palestinian,
årets	year,
efterhand	post,
piano	piano,
styras	controlled,steered,
drabbades	affected,where hit by,
julius	julius,
musikaliska	musical,
rådgivare	counsellor,advisor,
valla	wax,valla,herd,
jude	jew,
allvarlig	serious,
domkyrka	cathedral,abbey,
humle	hops,hop,
generell	general,
karibiska	caribbean,
musikaliskt	musical,musically,
anpassat	adapted,
uppväxt	growing up,
bönorna	bean,beans,
dokumenterade	documented,
utdelades	distributed,awarded,
hemligt	secret,
annorlunda	otherwise,
hemliga	secret,
främja	further,promote,promoting,
frivilligt	voluntarily,voluntary,
speglar	mirror,mirrors,
avrättning	execution,
frivilliga	volunteers,optional,
kina	china,
stöter	thrust,run,
simning	swimming,
regeln	rule,
muslimerna	muslims,the muslims,
inriktad	oriented,intent,
etablerat	established,
tvserien	the tv show,television program,
levt	survived,
fascism	fascism,
sydliga	southern,
familjens	the familys,family,
flög	fly,flew,
fenomen	phenomena,phenomenon,
leva	live,
utrikespolitiska	foreign policy,
väntan	awaiting,waiting,wait,
marknad	market,
kroniska	chronic,
beror	is,
stridande	conflict,
persons	a person's,persons,
japanska	japanese,
väntat	expected,
väntas	expected,
väntar	expect,
faser	phases,
orter	varieties,locations,
kartor	maps,
bushs	bush,
orten	resort,the suburb,
födelse	date,birth,
komplicerat	complex,complicated,
iberiska	iberian,
fasen	phase,
rapport	report,
fartyg	vessel,ship; vessel,
böcker	books,
kämpade	fought,
välja	select,
wallace	wallace,
undervisningen	teaching,the education,
sätt	manner,way,
organisation	organization,
behandlingen	the treatment,the treament,treatment,
spelarna	players,
klassen	the class,
tjänstemän	officers of,officals,officials,
marleys	marley's,marley,
passar	suitable,
hergé	herge,hergé,
femte	fifth,
märta	märta,
hamilton	hamilton,
karlsson	karlsson,
tredjedel	a third,third,
hotar	threatens,
term	term,
opera	opera,operator,
snabb	instant,
namn	name,
futharkens	futharkens,the futhark's,
viggo	viggo,
alternativ	alternative,
hotad	threatened,
färger	color,colors,
bildning	education,form,
semifinal	semifinals,semi finals,
förhandlingarna	negotiations,
stående	standing,above,
valuta	exchange,
rastafari	rastafarian,
amerikansk	american,u.s.,
åsikt	opinion,
tillhörighet	affiliation,belonging; affiliation,
behandlas	treated,
upprepade	repeated,
accepterad	acceptable,
stortorget	stortorget,the main square,
årliga	annual,
profil	profile,
accepterar	accepts,accept,
accepterat	accepted,
kent	kent,
variant	variant,variety,
juldagen	christmas day,
zuckerberg	zuckerberg,
etanol	ethanol,
nått	reached,
hjalmar	hjalmar,
gallien	gaul,
soundtrack	soundtrack,
arbetet	work,the work,
händelse	event,handel,
traditionen	the tradition,tradition,
motion	motion,exercise,
traditioner	traditions,
place	place,
någonsin	ever,
politiken	policy,the politics,
hemsida	homepage,
blood	blood,
origin	origin,
begår	commits,commit,
såldes	sold,
självbiografi	autobiography,selfbiografi,
centralamerika	central america,
george	george,
respekt	respect,
given	given,
nuvarande	current,
vågor	waves,
skjuten	shot,
cullen	cullen,
bahamas	bahamas,
skjuter	slide,
givet	granted,given,
hud	skin,
personlighetsstörningar	personality disorders,
spelats	recorded,been played,played,
webbplatser	webbsites,websites,
kronprinsessan	crown princess,
användandet	usage,use,
grund	because,
montenegro	montenegro,
alan	alan,
kallade	called,
hur	how,the,cage,
hus	house,a house,
webbplatsen	webpage,the website,site,
population	population,
smeknamn	nickname,
modellen	model,the model,
balans	balance,
marinen	navy,marines,
löfte	promise,
genomsnittet	average,the average,
framställning	preparation,production,
landsting	county,
modeller	models,
bildades	formed,was formed,
hjärtat	heart,the heart,
rena	pure,
mottagare	recipient,receiver,
ana	feel,ana,
anc	anc,
kromosomerna	chromosomes,the chromosomes,
maten	the food,
mando	command,
rent	clean,
jordskorpan	earth's crust,earth crust,
världen	world,the world,
avstånd	distance,
förste	the first,first,
första	first,
fysikaliska	physical,
förhållandena	conditions,the conditions,
gustavs	gustavs,gustav,
kust	coastal,coast,
periodvis	periodically,
stjärnornas	stellar,the star's,
knutna	associated,attached,tied,
diskussioner	discussions,discussion,
falla	fall,
 miljoner	one million,millions,millon,
invånarna	inhabitatants; citizens',residents,
staterna	usa,
täckt	covered,
täcks	covers,
lisbet	lisbet,
astronomiska	astronomical,
erkänner	admits,recognize,
stövare	beagle,hound,
täcka	cover,thank,
tron	faith,
ronaldinho	ronaldinho,
mänskligheten	humanity,
bernadotte	bernadotte,
isolering	isolation,
tros	belived,
tror	believe,think,
bandets	the bands,band,
gula	yellow,
tvprogram	tv program,tv-show,
guld	gold,
tidningarna	papers,
flydde	fled,
motivet	the motive,subject,
ovanligt	unusual,
gult	yellow,
iväg	away,off,
ovanliga	unusual,rare,
analys	analysis,
berättelser	stories,
webbkällor	web sources,
larsson	larsson,
aktiviteten	activity,
grundandet	founding,
tränaren	coach,
jazz	jazz,
administrativ	administrative,administration,
nedåt	down,down; downwards,
väder	weather,
ansågs	was,seemed,
forsberg	forsberg,
beredd	prepared,
tränade	trained,
dramat	drama,the drama,
umeå	umeå,
joker	joker,
republika	republic,
osäkert	insecure,unclear,uncertain,
baltikum	the baltics,baltics,
förmån	benefit,advantage; in favor of; benefit,
minnen	memories,memory,
underlätta	ease,facilitate,
tekniska	technical,
inspelningen	recording,
uppdraget	task; assignment,assignment,
tekniskt	technical,
college	college,
stanley	stanley,
minnet	memory,
älg	elk,moose,
freden	the peace,peace,
federal	federal,
utbud	availibility,
skett	done,happened,
önskade	desired,wished,
hämtar	download,is,
återigen	once again,yet again,aterigen,
intresserad	interested,
hämtat	collected,taken,
konstnären	artists,the artist,artist,
mellan	between,
antagligen	probably,
konstnärer	artists,
bekämpa	combat; fight,fight,
ruiner	ruins,
dödade	killed,
myter	myths,
högre	higher,
come	come,
summa	sum,total,
sydeuropa	southern europe,
region	region,
ordagrant	literal,verbatim,
spindlar	spiders,
lenins	lenin,lenin's,
introducerades	introduced,
gjorde	did,
gjorda	made,done,
pakistan	pakistan,
utgåvor	editions,issues,
regler	rules,
period	period,
pop	pop,
fransk	french,france,
werner	werner,
statens	state,the government's,
utformning	layout,formation,
hävda	claim,asserting,
poe	poe,
skånska	scanian dialect,scanian,
howard	howard,
folken	the peoples,people,
strikta	strict,
förekomsten	existence,presence,
dagarna	the days,day,
musikstil	music,music style,
folket	the people,people,
invaderade	invaded,
anderna	andes,the andes,
sändebud	envoy,
andres	andres,other's,
stadshus	city hall; town hall,town hall,
tjänster	services,
kapitulation	surrender,capitulation,
tiger	tiger,silent,
övrig	other,
minister	minister,
epok	epoch,
kaos	chaos,
champions	champions,
hughes	hughes,
användes	was used,
riktade	targeted,
bilderna	the pictures,
influenser	influence,influences,
cash	cash,
arnold	arnold,
spreds	spread,
ifrån	off,
fiende	enemy,
grundlagen	constitution,the constitutional law,
odens	odin's,node,oden's,
universums	universe,universe's,
pippi	birdie,pippi,
hamn	harbor,port,
nyare	newer,
knyta	tie,
grönland	greenland,
status	status,
producera	produce,producing,
republikens	republic's,republic,
fysiologi	physiology,
protoner	protons,
hjärta	heart,
linjerna	the lines,lines,
göring	goring,cleaning,
privilegier	privileges,
vatikanstaten	vatican city,vatican,
relaterade	related,
modet	courage,fashion,
medvetna	aware,conscious,
kommunistisk	communistic,communist,
breda	wide,
hårdvara	hardware,
without	without,
tjänsten	service,
nordkoreas	north korea,north coreas,
medellivslängd	average lifespan,life expectancy,
arkitekten	architect,the architect,
kopplingen	coupling,
lyckan	happiness,
fördelas	distribute,distributed,
listorna	menus,the lists,
kommentarer	comments,
förklarades	was explained,explained,
ekologiska	ecological,
enligt	according (to),according to,
kill	kill,
knäppupp	knäppup,knäppupp,
harrison	harrison,
moçambique	mozambique,
leta	search,check,
utvinns	extracted,
starka	strong,
tim	tim,h,
rose	rose,
regent	regent,
rosa	pink,
utbyte	yield,trade,
starkt	strongly,strong,
lett	resulted,
utvinna	extract,
pendeltåg	commuter,
delstat	state,land,
guldbollen	golden ball,guldbollen,
ross	ross,
riket	kingdom,the land,
mesta	most,
porto	postage,
vampyren	the vampire,vampire,
delhi	delhi,
utrikespolitik	foreign policy,foreign affairs,
uppslagsordet	lookup word,lexical entry; word,
kille	guy,
tid	time,
majoritet	majority,
inflation	inflation,
vampyrer	vampires,
walk	walk,
riken	the kingdoms,kingdoms,
kommentar	comment,
afrikas	africas,africa,
talrika	numerous,
mexikanska	mexican,
cooper	cooper,
anföll	attacked,
rammstein	rammstein,
verksamheten	activity,
madrid	madrid,
styrkor	strenghts,forces,
teorin	theory,the theory,
gång	once,time,
passera	pass,
latinet	latin,
alkoholer	alcohols,
verksamheter	operations,businesses,activity,
försvarare	defenders,defender,
tiders	days',times,
fiktion	fiction,
inspirerades	inspired,
sitta	sit,
stopp	stop,
moon	moon,
härledas	derived,
lärda	scholars,savants,
buddha	buddha,
lärde	learned,
uppbyggnad	construction,
publicerat	published,
storhetstid	heyday,
liberala	liberal,
football	football,
servrar	servers,
geografi	geography,
genom	through,
tyskt	german,
korrekt	correct,
mandelas	mandelas,mandela's,
tyska	german,
tyske	german,
förbindelser	relations,
on	on,
om	of,if,
indianska	red indian,native american,
spelet	the game,game,
og	og,
of	of,av,
oc	o.c.,oc,
stand	stand,
nåddes	reached,
os	os,
spelen	the games,
befäl	command,
koppling	clutch,connection,
cambridge	cambridge,
ansträngningar	effort,
tolkning	interpretations,
domstol	court,
överföras	transfer,transferred,
befinna	be,
mental	mental,
medlemsstaternas	member,member state,
fisk	fish,
valley	valley,
serbien	serbia,
förrän	until,
jul	christmas,
inriktning	direction,orientation,
uppåt	up,upwards,
ingredienser	ingredient,ingredients,
manuskript	manuscript,script,
varning	warning,
ämbetsmän	officer,bailies,officers,
chaplin	chaplin,
kvinnornas	womens,women,
taylor	taylor,
felix	felix,
närmast	nearest,closest,mediately,
fjorton	fourteen,
pengar	money,
ökning	increase,
operation	operation,
köpenhamn	copenhagen,
många	many,
roses	roses,
mötley	mötley,
utgifter	expenditure,expenses,
babylon	babylonia,babylon,
visade	showed,showed; displayed,
separata	separate,
grupp	group,
sällskapet	society,the company,
symbol	symbol,
erövring	conquest,
missbruk	abuse,
vinnaren	winner,
observatörer	observers,
symtomen	symptoms,ymptoms,
villkor	conditions,
distriktet	district,
barcelona	barcelona,
calle	calle,
erfarenhet	experience,
visby	visby,
all	any,
ali	ali,
alf	alf,
separat	seperate,separate,
samhället	the society,society,
stödde	supported,
samhällen	communities,societies,
utomliggande	external; ex-territorial,outlying,
sakrament	sacrament,
antogs	adoption,was assumed,
uppdrag	job,missions,
persiska	persian,
funktionerna	functions,the functions,
brottet	offense,the crime; offense; infraction; transgression,
röstade	voted,
ögonen	eyes,
gary	gary,
påstående	claim,assumption,
program	application,
cykeln	cycle,
kvar	left,
löper	runs,at,
färgerna	colors,
liter	liters,
litet	small,
oavgjort	tie,draw,
song	song,
far	father,
fas	phase,
fat	barrel,
runtom	throughout,around,
simpsons	simpsons,
fan	devil,fan,
sony	sony,
liten	small,
unionens	the union,the union's,
tjeckiska	czech,
choklad	chocolate,
knutsson	knutsson,
list	cunning,
kopplas	connected,coupled,
förtryck	opression,
lisa	lisa,
över	over,
iran	iran,
hitta	see,come up, find,
grekland	greece,
ted	ted,
istiden	ice age,the ice age,
tex	for example,e.g.,
design	design,
haag	the hague,
what	what,
enklaste	easiest,
sun	sun,
vaginalt	vaginal,
kinesiska	chinese,
version	version,
spelning	gig,playing,
sur	sour,
mördades	murdered,was murdered,
guns	guns,
fäste	bracket,
christian	christian,
dottern	the daughter,daughter,
upptäcka	discover,
regerade	reigned,
avrättades	was executed,executed,
leeds	leeds,
madeleine	madeleine,
upptäckt	discovered,found,discovery,
norden	scandinavia; (nordic area; region),the nordic countries,north,
nordens	the scandinavian countries',scandinavia,nordic,
upptäcks	discoverd,detected,is discovered,
råder	advises,is,
kommande	upcoming,
soloalbum	solo album,
kärnvapen	nuclear,nuclear weapons,
tillhörde	belonged to,belonging to,
magnitud	magnitude,
arabemiraten	united arab emirates,uae,the arab emirate,
nyfödda	newborn,
snus	snuff,
uppkomst	origin,onset,
kategorispelare	category player,
filmerna	films,the movies,
stöd	support,
syfte	purpose,
syfta	aim,refer,
smak	taste,flavoring,
socialdemokraterna	members of the social democracy,social democratic,
anarkism	anarchism,
succé	succession,
kommittén	the committee,committee,
branden	the fire,
förebild	role model,
autonom	independent,autonomic,
bekräftade	confirmed,
genomsnittliga	average,
israel	israel,israeli,
permanenta	permanent,
alltid	always,
akademiens	academy,the academy's,
glas	glass,
hålet	hole; gap,hole,the hole,
floyd	floyd,
glad	happy,
östra	eastern,
naturligt	natural,
legender	legends,
godkänt	approved,pass,
decenniet	decade,
decennier	decades,
kryddor	spices,
förhåller	relate,relationship,
naturliga	natural,
pony	pony,
duett	duet,
bosatt	resident,lived,
styrs	is controlled,ruled,
elektrisk	electric,elektirsk,
historiskt	historic,historically,historical,
court	court,
breaking	breakingpoint,breaking,
brittisk	british,
satanism	satanism,satanic,
historiska	historical,
härstamning	lineage,origin,descent,
välgörenhet	charity,
indelade	divided into,
rocksångare	rock singers,rock singer,
taget	a time (practically; virtually; any; at all),time,
sven	sven,
tagen	taken,
grundämne	elemental,element,
fötterna	feet,
ångest	anxiety,
fötts	born,borned,
atomer	atoms,
regnar	rains,raining,
anarkistiska	anarchist,
praktiska	practical,
bildade	formed,
tsar	tsar,czar,
homosexuella	homosexual,gay,
grande	grande,grand,
greklands	greek country,
människors	humans,human,
friidrott	athletics,track and field,
längs	along,
avvisade	rejected,
september	september,
sträckte	extended,
emmanuel	emmanuel,
mission	mission,
australien	australia,
längd	length,
retoriska	rhetorical,
hounds	hounds,
islam	islam,
lyder	reads,obeys,
rika	rich,
abbey	abbey,
centralort	central city,centralot,
rikt	target,rich,
stadsparken	city park,
prag	prague,
stephen	stephen,
argentina	argentina,
jämte	plus,
fenomenet	the phenomenon,phenomenon,
kategorieuropeiska	european category,
styret	gate,
medborgerliga	civil,
kärna	core,quarks,
postumt	posthumously,
landborgen	the ridge,
marcus	marcus,
försöken	attempts,the tries,
journalisten	journalist,the journalist,
forna	former,
stilen	style,
slidan	vagina,vaginal,
journalister	journalists,
försöker	try,tries,trying,
principer	principals,principles,
kustlinje	coastline,
ringar	rings,
drycken	the drink,
betyg	grades,
hawaii	hawaii,
konstnärlig	art,artistic,
aldrig	never,
drycker	beverages,
stenar	stones,blocks,
ollonet	penis head,glans,the glans,
därvid	thus; thusly; then,therewith,
nepal	nepal,
europas	europe,
hill	hill,
väg	vague,way,
kvinna	woman,
väl	selecting,good,
vän	friend,
helgdagar	holidays,
poliser	police (-men; -women),police,
ökad	increase,increased,
islamistiska	islamist,
densiteten	density,
beräknades	calculated,estimated,
ökat	increased,
spelades	filmed,
kritiserar	criticize,
polisen	police,
faller	fall,
fallet	case,the case,
stavningen	the spelling,
konsumtionen	consumption,
fallen	case,cases,
aminosyror	amino acids,
filosofins	philosophy,the philosophy,
heinz	heinz,
colombia	colombia,
pablo	pablo,
bland	inter,including,
blanc	blanc,
story	story,
infört	introduced,
lördagen	the saturday,saturday,
automobile	automobile,
misslyckas	fail,fails,
harris	harris,
stort	large,big,
motiveringen	the motivation,ground,
storm	storm,
kristendomens	christianity's,christianity,
brasiliens	brazil's,
ecuador	ecuador,
familjerna	families,
mikael	mikael,
gränser	borders,frontiers,
hotel	hotel,
kongress	congress,
serotonin	serotonin,
framtiden	future,the future,
hotet	the threat,threat,
fattigaste	the poorest,
gränsen	limit,border,
besökare	visitors,
siffra	number,figure,
king	king,
illegala	illegal,irregular,
matcherna	the games,
direkt	direct,directly,
nöd	distress,emergency,
pjäsen	play,piece,
dans	dance,
kategorisommarvärdar	category summer hosts,
guden	god,the god,
stjärnan	star,the star,
tillåta	allowing,
klubb	club,
anläggningar	plants,facilities,
kusin	cousin,
tilldelas	assigned,
tabell	table,
omskärelse	circumcision,
slåss	fight,
divisionen	division,
wilson	wilson,
väsen	being,
bedriver	conducts,operate,
inriktningar	specializations,
unga	young,
jämförelsevis	comparative,in comparison,comparatively,
judas	judas,
judar	jews,
kiss	view,
folkgrupper	communities,ethnic groups,
electric	electic,electric,
dagliga	daily,
park	park,
stjärnans	star's,the stars,
dagligt	daily,
industrialiserade	industrialized,
agnostiker	agnostic,agnostics,
sånger	songs,
mineral	minerals,mineral,
windows	windows,
salt	salt,
influensan	the influenza,flu,
sången	the song,song,
borgmästare	mayor,
statsskick	polity,form of government,government,
kosovo	kosovo,
tjugo	twenty,
ursprungliga	original,
kapitulerade	surrendered,
tilly	tilly,
månen	the moon,man,
tills	until the,until,
beräkningar	calculations,
canaria	canaria,
bidrog	contributed,
moses	moses,
hit	to here,here,
hiv	hiv,
stormakterna	great powers,
inklusive	including,
vardera	either,each,
fattiga	poor,
jobbade	worked,
händer	happening,hands,
sofie	sofie,
solsystemet	the solar system,
utvidgade	expanded,
tvkanaler	tv channels,
mediciner	medicines,
knapp	button,bare,
tidszon	timezone,time zone,
vincent	vincent,
norrköping	norrköping,
poäng	score,
virginia	virginia,
utsatt	exposed,
bars	bar,
etiopien	ethiopia,
art	kind,art,
bart	offense,bart,
arv	heritage,
fiske	fishing,
bara	only,
are	are,
arg	angry,
flyttade	moved,
stjäla	steal,
arm	arm,
barn	child,
pär	pär,
bortsett	except,
planeras	is planned,planned,
planerar	plan,planned,
uppskatta	appreciate,
inga	not,no,
planerat	planned,
invaldes	was elected,
planerad	planned,
muslim	muslim,
verksamhet	work,activity,
där	where,in which,
intäkter	revenues,incomes,
herrar	gentlemen,men,
uppkom	arose,
godkändes	approved,
tiderna	the times,times, ages,time,
balkanhalvön	balkan peninsula,
startades	started,
operan	opera,
roman	novel,
lägret	the camp,camp,
påstår	states,claims,asserts,
hypotesen	the hypothesis,
lära	lara,get to know,learn,
borta	gone,
vidare	moreover,furthermore,
lärt	learned,learnt,
stärktes	was strengthened,strengthened,was strenghten,
belägna	located,disposed,
besegrade	defeated,
östtyskland	east germany,
utifrån	from,
hypoteser	hypotheses,hypothesis,
ps	ps,p.s,p.s.,
java	java,
göteborg	gothenburg,
personalen	personnel,the staff,
kungafamiljen	the royal family,
johannes	johannes,john,
avslutade	ended,finished,
byxor	pants,
resultat	results,result,
ph	ph,
pi	pi,
chandler	chandler,
flight	flights,flight,
togs	taken,were taken,
publiken	audience,
sydafrikas	south african,south africa's,
rättigheterna	the rights,
gården	farm,courtyard; house; farm (-house),
konflikter	conflicts,conflict,
konflikten	the conflict,conflict,
deltog	participated,
sådan	such,
inspelningar	recordings,
ägs	is owned,owned,
styr	controls,
ris	rice,
rik	rish,rich,
sjöarna	the lakes,lakes,
byggnaderna	building,buildings,the buildings,
skeppen	the ships,
fysisk	natural,physical,
demografi	demographics,demography,
tidpunkten	the time,the moment,time,
ideologier	ideologies,
sjunkit	decreased,
förföljelse	persecution,
torbjörn	torbjörn,torbjorn,
spears	spears,
låtit	let,had,
bröllopet	the wedding,wedding,
byar	villages,
skåne	skåne,
uppbyggd	structered,structured,built-up,
författare	author,
uppbyggt	structured,
kokpunkt	boiling point,
vinklar	angle,angles,
finansiera	fund,finance,
italiensk	italian,
sjunga	access,sing,
höjer	raising,
edge	edge,
vetenskapen	the science,science,
kyrkans	the church's,church,
alfabet	alphabets,alphabet,
uttalande	statement,
kontinentala	continental,
komplett	complete,
konstitution	constitution,
påverkade	influenced,
remmer	remmer,
dåtidens	past times,that time,
prince	prince,
namnet	name,
folkräkning	census,
skalv	quake,
minoriteter	minorities,
bostad	lodge,property,
omedelbar	instant,immediate,
försvunnit	disappeared,
skall	is,shall,
minoriteten	minority,
idé	ide,
emigrerade	emigrated,
px|centrerad	px | centric,
skala	scale; size,scale,
färdiga	finished,
synnerhet	specially,particular,
djupare	depth,deeper,
rastafarianerna	rest are faria,
begravdes	buried,
användas	used,
stoppade	stop,stopped,
upplevelse	experience,
exakt	accurately,
våldsamma	violent,
näringsliv	business,
banbrytande	groundbreaking,
sammansättning	composition,
hittar	found,finds,
hittas	found,
hittat	found,
minskning	decline,
landskommun	rural municipality,
norrut	north,
sjöfart	sea voyage,maritime,
kongo	congo,kongo,
lettland	latvia,
trummis	drummer,
global	global,
förteckning	listing,
flottan	the fleet,navy,the navy,
thailand	thailand,
huvudstad	capital,
låtarna	the songs,songs,
ungefär	approx.; approximately,about,
höjden	height,
föräldrar	parents,
grekerna	greek,greeks,
prov	test,
frälsning	salvation,
fungera	act,
anne	anne,
trinidad	trinidad,
höjdes	increased,was raised,
höjder	altitudes,heights,
turism	tourism,
diamant	diamond,
palmes	palme,plame's,
ställningen	position,
tävlade	competed,
presenteras	presented,
anklagades	accused,
judendom	judaism,jewism,
kostnaderna	costs,the costs,
grundläggande	because lag of,primary,fundamental,
påtryckningar	pressures,pressure,
tätt	tight,tightly,
virus	virus,
ande	of,spirit,
dialog	dialogue,
täta	close,seal,
socialistisk	socialistic,socialist,
oktoberrevolutionen	the october revolution,october revolution,
genomföras	carried out,be performed,
medborgarna	the citizens,citizens,
reglerna	rules,rules; regulations,
hållet	cohesive,way,
abbas	abbas,
km²	square kilometre,
laget	the team,stroke,
håller	is,holds,
dricka	drinking,drink,
fast	solid,though; although; fixed; permanent,even though,
jugoslavien	yugoslavia,
bagge	bagge,
bruk	using,use,
laila	laila,
ateister	steister,
delning	pitch,
rasade	collapsed,
regionen	the region,region,
längtan	longing,
sköter	handles,handle,
kritikerna	critics,the critics,
delta	participate,delta,
tidigast	the earliest,
junior	junior,
medeltidens	ages,medieval,
anklagelser	allegations,
planeternas	the planets,planets,the planets',
världskrigen	the world wars,world wars,
styrande	rulers,governing,
aktier	share,
världskriget	world war,
guyana	guyana (name),guyana,
tolka	interpreting,interpret,
handels	commercial,
z	z,
tidens	time's,
svenskspråkiga	swedish speaking,
ägdes	owned,
singlarna	singles,
tidpunkt	date,time,
home	home,
däribland	including,
graham	graham,
veckorna	weeks,
rainbow	rainbow,
stadion	stadium,
möten	meetings,
höga	high,
psykoterapi	psychotherapy,
högst	highest,maximum,
mötet	the meeting,meeting,
hanen	the cock,male,
urval	selection,
skyddas	protected,(is/are) protected,
skyddar	protection,protects,
sutra	sutra,
beräknas	calculated,
beräknar	computes,values,
tittarna	the viewers,viewers,
medina	medina,
stadigt	stable,steadily,
konvertera	convert,conversion,
betyder	means,
råkar	happens,happens to,
jugoslaviska	yugoslav,yugoslavian,
modernismen	modernism,
klubbens	club,
oväntat	unexpected,
underlättar	facilitates,
vice	vice,
europeiska	european,
parallella	parallel,
microsoft	microsoft,
nasa	nasa,
karma	karma,
lagstiftning	law-making,regulation,
europeiskt	european,
nash	nash,
förhandla	negotiate,negotiating,
psykologi	psychology,
beträffande	on,
kanal	channel,
steve	steve,
jimi	jimi,
stieg	stieg,
moseboken	genesis,
kolonialismen	the colonialism,colonialism,
simon	simon,
uppmaning	call; injunction,call,exhortation,
fortfarande	still,
romerna	the romani,the romani people,
kazakstan	kazakstan,
generellt	generally,
generella	overall,general,
hinduism	hinduism,
fotnoter	footnotes,
pengarna	the money,money,
varierar	varies,vary,
vapen	weapons,weapon,
kategoritvseriestarter	category television series starts,
varierat	varied,
mesopotamien	mesopotamia,
sjukdomar	diseases,disease,
medverkade	participated; contributed,participated,
kommitté	committee,
avslutas	close,ends,closing,
avslutat	completed,
tvinga	force,
historikern	historian,
demokratiskt	democratic,
äta	eat,
inleder	start,initiates,
noter	notes,notation,
öron	ear,
läkemedel	medicine,
utanför	outside,
melodier	melodies,
byggd	built,
reptiler	reptiles,
bygga	building,build,
indirekt	indirectly,
skadad	damaged,
åtminstone	at least,
århundradet	century,
skadan	damage,
influerad	influenced,
anderssons	anderssons,andersson's,
skadas	damaged,
västlig	western,
konstant	constant,
folk	public,people,
influerat	influenced,
hölls	was held,was,
assisterande	assistant,assisted,
kris	crisis,
skrivna	written,
judy	judy,
krig	war,
dramatiska	dramatic,
bröts	was fractured,broke,
insats	stake,
koloni	colony,
hdmi	hdmi,
producenten	the producer,producer,
turismen	tourism,
producenter	producers,
diamanter	diamonds,
åtgärder	measures,
filosofi	philosophy,
astrid	astrid,
tvingats	forced,had,
fauna	fauna,
buddhistiska	buddhistic,buddhist,
ukraina	ukraine,
metro	metro,
innehar	holds,
innehas	held,occupied,
innehav	owning,
springsteens	springsteen's,springsteens,
plattan	plate,
fortsätter	continues,continue,
populärkulturen	popular culture,
översättningar	translations,
tjänar	earns,serves,
zlatan	zlatan,
reda	out,find our,
gemenskap	fellowship,community,
föreställande	depicting,
motor	engine,
juryns	the jury's,jury,
redo	prepared,
varpå	thereafter,whereupon,
from	from,
bestämmelser	measures,conditions,
usa	united states of america,usa,
fel	errors,error,
fem	five,
sevärdheter	attractions,
upplöstes	dissolved,
källorna	source,the sources,
inlandet	inland,the inland,
öppnat	opening,
andliga	spiritual,
penis	penis,
införande	introduction,
hindrade	prevented,
vägrade	refused,
fungerar	works,
reguljära	regular,
beskriva	describe,
automatiskt	automatic,
beskrivs	described,
tar	takes,
tas	is,is taken,
föreslår	suggests,suggest,
platser	points,places,
crick	cricket,crick,
engels	engels,
treenigheten	tinity,the trinity,trinity,
tag	while,
hilton	hilton,
tal	speech,
kanadensiska	canadian,
sir	sir,
ondska	evil,
löften	promises,
notation	notation,
six	six,
brian	brian,
sig	to,itself,
undantaget	except,
sin	its,
väpnad	armed,
kostym	costume,
kontroversiellt	controversial,
förekommande	occuring,where,
oavsett	whether,regardless; whether; irrespective of,regardless,
tack	thanks,
religiös	religious,
bertil	bertil,
kategoriwikipediabasartiklar	category wikipedia basartiklar,
kontroversiella	controversial,
eritrea	eritrea,
light	light,
centralorter	centers,
framförts	forward,
öresund	Øresund,the sound,
jolie	jolie,jolies,
besegrat	defeated,
mekka	mecca,
blandad	mixed,blended,
skapande	building,creative,
företrädare	representatives,
elin	elin,electrical,
förklaras	explained,
elit	elite,
blandat	mixed,
karlstad	karlstad,phoenix,
blandas	mixed,mixes,
spotify	spotify,
stiga	rise,rising,
uppmärksammad	noted, come to attention,attention,noticed,
terriers	terriers,
befolkning	population,
byn	village,
floder	rivers,
permanent	permanent,
försvar	defence,defense,
lärjungar	disciple,
thåström	thåström,thastrom,
carola	carola,
skede	period,analysis,
cypern	cyprus,
verkligen	real,
washington	washington,
fler	more,
andlig	spiritual,
östtimor	east timor,
satelliter	satellite,
exempelvis	e.g.,
komma	access,
ale	ale,
billy	billy,
växande	growing,
konungariket	kingdom,
mätt	dull,
studios	studios,the studio's,
australiska	australian,
säsonger	seasons,
barnets	the childs,child,
byter	changes,exchanges,
kvarteret	quarter,the neighborhood,
säsongen	season,
studion	studio,the studio,
kritik	criticism,critisism,critique; criticism,
alger	algaes,algae,
förbjuda	ban,prohibiting,
uggla	owl,
minskad	decreased,reduced,
hantverkare	handy worker,craftsman,
fiktiva	fictitious,
svar	answer,response,
bål	prom,
nobelpristagare	nobel laureate (-s); nobel prize winner (-s),nobel laureates,
minskat	decreased,reduced,has decreased,
uppnå	achieving,achieve,
minskar	decrease,
förutsättningar	prerequisites,(pre-)conditions,condition,
hörs	heard,
hört	heard,heared,
hjälpt	helped,
vulkanutbrott	vulcano eruption,volcanic eruption,
utmärker	characterized,
höra	know,
hjälpa	helping,
york	york,
studioalbumet	studio album,
philip	philip,
domare	judge,
hörn	corner,
fotbollslandslag	football team,national football team,
gångna	past,past; gone,
anslutning	connection,
tyst	quiet,silent,
waterloo	waterloo,
barns	child,childrens,children,
via	through,
adrian	adrian,
tvserier	tv shows,tv-series,
tysk	german,
rudolf	rudolph,rudolf,
ovanpå	top,on top of,
revolutionens	revolution,the revolutions,
isbn	isbn,
brasilien	brazil,
velat	wanted,
nietzsches	nietzsche,nietzsche's,
värsta	worst,
regenter	monarchs,regents,
skyddade	protected,
nätverk	network,
enkelt	easy,
förhöjd	enhanced,elevated,
fågelhundar	bird dogs,
meddelanden	messages,
omfattning	extent,
misslyckande	failure,
sankta	sankta,saint,
diskutera	discussed,discuss,
rösträtt	vote,right to vote,
valde	selected,chose,
valda	chosen,
vingar	wings,
juli	july,
vind	wind,
dödligheten	mortality,
resterande	remainder,remaining,
belgien	belgium,
franska	french,
holland	holland,
franske	the french,french,
birgitta	birgitta,
tommy	tommy,
framgång	success,
algeriet	algeria,
franskt	french,
tomma	empty,
tyskarna	germans,the germans,
heydrich	heydrich,
fyrtio	forty,
cohen	cohen - it's a name,cohen,
benny	benny,
avgörs	determined,is determined,decided,
blir	become,is,
farligt	dangerous,hazardly,
ringen	ring,
gäng	group,thread,
intervju	interview,
storbritannien	great britain,uk,
byggas	prevented,build,
uppfann	invented,
lopp	course, passage,race,
ansåg	thought,found,considered,
besittning	dominion,possess,
kristi	kristi,
betydligt	considerably,
centra	center,
ström	power,
centre	centre,
who	who,
intogs	was taken,was captured,
representation	representation,
staternas	states,
öken	desert,
planerade	planned,
förbundsrepubliken	the federal republic,federal republic of,
undersökte	investigated,
regeringschef	head of government,government,
miljontals	millions,
enbart	only,
judendomen	judaism,
kategoriamerikanska	u.s. category,
moberg	moberg,
uefa	uefa,
blandade	mixed,
funktionella	functional,
debatt	debate,
julafton	chistmas eve,christmas eve,
pastoral	pastoral,
angående	concerning,reference,
dödades	were killed,killed,
asterix	asterix,
rösten	rust,the voice,
nilsson	nilsson,
filmer	films,movies,
röster	votes,
beroende	dependent,
hållning	position,entertainment,
allmänhet	in general,general,
träffa	meet,see,
gränsar	adjacent,
heta	hot,be named; be called,be called,
överens	in agreement,
gudar	gods,
linje	line,
presley	presley,
hett	hot,
närstående	relative,relatives,kindred,
samtycke	consent,
städer	urban,cities,
begäran	request,
förbinder	connects,undertake,
torka	dry,
respektive	and,respective,
mestadels	mostly,
kvinnorna	the women,women,
berömd	famous,
nationernas	the nations,nations,
rikare	richer,
motståndare	opponents,opponent,
theta	theta,
funktion	function,
upplysning	enlightenment,
praktisk	practical,
sydstaterna	southern states,southern united states,
faktiskt	in fact; actually; indeed,really,actually,
vandrar	wanders,migrates,
joe	joe,
swift	swift,
jon	jon,
sångaren	singer,the singer,
allsvenskan	headlines,
ingemar	ingemar,
påtagligt	substantially,considerably,markedly,
utvecklingen	development,the development,
teoretiker	theorists,
kolhydrater	carbohydrates,
april	april,
västerländsk	western,
brons	bronze,
vattnets	water,the water's,the waters,
bronx	the bronx,
förespråkare	spokesman,proponent,
betecknar	represent,denotes,represents,
betecknas	labelled,denote,
kategorityska	category: german,
exakta	exact,
korruption	corruption,
wall	wall,
vittne	witness,
publicerad	published,
walt	walt,
cirka	about,approximately,
utsedd	appointed,
innebära	mean,
publiceras	publishes,published,
framträdanden	appearances,
jenny	jenny,
utkom	issued,
klara	clear,
dödshjälp	euthanasy,euthanasia,
hindu	hindu,
kopplade	connected,
bbc	bbc,
beskrivning	description,
månar	moons,
klart	clear,done,
månad	month,
strindbergs	strindberg's,strindberg,
ständig	constant,
naturtillgångar	natural resources,
mike	micke,mike,
liverpool	liverpool,
nickel	nickel,
väljs	selected,
turneringen	the tournament,
dominera	dominate,
lutherska	lutheran,
försvann	disappeared,
hms	hms,
fortsättningen	the continuation,remain,
neutrala	neutral,
deklarerade	declared,
last	load,
plikter	duties,
present	gift,
godkännande	approval,authorization,
bråk	brawl; fight,fights,fraction,
problemen	problems,the problems,
officiell	official,authentic,
största	biggest,maximum,largest,
anpassa	adjust,
will	will,
fördelade	divided,distributed,
nominerades	was nominated,nominated,
wild	wild,
fjärdedel	quarter,fourth,
folktro	popular belief,folklore,
explosionen	the explosion,
sagan	story,
vuxit	grown,
gemensamt	single,in common,
bosättare	settlers,
syftar	refers,seek to,
motiv	subjects,motif,
jehovas	jehovas,jehova's,
röra	move,
uppstå	develop,occur,
ramels	ramel's,
varar	duration,lasts,
buddhism	buddhism,
pojkar	boys,
samband	connection,
inch	inches,
skickade	sent,
gett	given,gave,
annekterade	annexed,annexation,
tvister	conflicts,disputes,
mottagande	host,reception,
övervägande	predominant,predominantly,
romeo	romeo,
romer	romani people,roma,
student	student,
raka	straight,
rätt	right,entitled,
misstag	error,mistake,
klubbar	clubs,
vilar	rests,
banden	bands,bander,the bound,
terrorismen	terrorism,the terrorism,
undersökningar	surveys; investigations,studies,
moderaterna	the moderates,moderates,
ekosystem	ecosystem,eco system,
övertyga	convince,
english	english,
bandet	band,
organisationens	organization,the organizations,
hårdrocken	hard rock,
lön	salary,wage; salary,
biologisk	biological,
singeln	single,
mfl	etc,etc.,
möjligheter	potential,
uppkommer	arises,arises; generated,
möjligheten	the ability,
rachels	rachel's,
erfarenheter	experiences,experience,
högskolor	colleges,
förtroende	confidence,
miljöer	environment,environments,
antisemitism	antisemitism,
rocken	rock,
brutit	cut; break,broken,
mytologiska	mythological,
jarl	earl,jarl,
genombrottet	break-through,breakthrough,
alldeles	completely,altogether,
hoppa	skip,drop out,
bell	bell,
sky	sky,
rättsliga	justice,legal,
engelsk	english,
ske	be,happen,
ska	will,
fyller	turns,turn; fill,
sanskrit	sanskrit,
hotade	threatened,
psykoser	psychoses,
färgen	color,the color,
olle	olle,
agerande	behavior,
älska	love,
know	know,
press	press,
psykosen	psychosis,the psychosis,
säljs	sold,
georges	georges,
budet	the bid,the commandment,
miami	miami,
djupa	deep,
huruvida	whether,
sälja	sell,
gorbatjov	gorbachev,
immunförsvar	immune defense,
finansieras	financed,funded,
djupt	deep,
säkra	reliable,safe,secure,
serbiska	serbian,
tjeckoslovakien	czechoslovakia,
handeln	trade; commerce,trade,
berömt	famous,praised,
bibliska	biblican,biblical,
efterfrågan	demand,
gäst	guest,
export	export,
försvinna	vanish,
star	star,
skandinavien	scandinavia,
använts	was used,used,
genomsnitt	average,
planering	planning,
trianglar	traingles,
gammalt	old,
risker	risker,
undviker	avoid,
klassificera	classifying,classify,
setts	observed,seen,
mankell	mankell,
låter	let,
låten	the song,song,
sjunker	flag,sinks,
markera	mark,
utsöndras	exudes,secreted,
uppvärmning	heating,warming,
mitt	my,center,
slut	end,out,
dateras	dates,dated,
sommarspelen	summer games,summer olympics,
lång	long,
ljung	heather,
låna	borrow,lana,
pressfrihetsindex	press freedom index,
substantiv	noun,
tillräcklig	sufficient,enough,
överlevde	survived,
bestämma	determining,decide,
oberoende	independent,
avsnittet	episode,
saken	the thing,matter,
saker	things,items,
avsnitten	sections,chapters,
mäta	compare,feeding,
främre	forward,front,
egna	own,
återvänt	returned,returning,
någorlunda	fairly,somewhat,
avrättade	executed,
tillbringade	spent,
mäts	is measured,
sektorn	sector,the sector,
floden	river,the river,
vidta	take,
flyger	flies,flying,
stressorer	stressors,
glukos	glucose,
folkpartiet	liberal party,
konstruktion	construction,structure,
födelsetal	birthrate,birth rate,
citat	quote,
val	choice,
idén	the idea,idea,
vad	as,
smeknamnet	nickname,
mäter	measuring,measure,
var	was,
regisserad	produced,directed,
vacker	beautiful,
nordamerikanska	north american,
lundell	lundell,
granne	neighbor,
hundratal	hundred,
ingått	entered,entered into,
krigsslutet	end of war; war's end,
stadens	the town's,the citys,city's,
karta	map,maps,
made	made,
rybak	rybak,
arne	arne,
tema	theme,
missnöjet	grievance,discontent,
kuriosa	curiosities,trivia,
reaktorn	reactor,
problemet	the problem,
stormakter	world powers,great power,superpowers,
eu	eu,
utöva	carry,exercise,
runor	runes,
kant	kant,
året	the year,all year,years,
illinois	illinois,
book	book,
ursprunget	origin,
åren	the years,years,
intresse	interest,
juni	june,
behandlar	treats,treat,
tolkas	is interpreted,interpretation,interpret,
tolkar	interprets,
shakespeares	shakespeare's,shakespeare,
tvfilm	tv movie,
personligen	individual,personally,
fira	celebrate,
ställningar	positions,notions,
margaret	margaret,
markant	considerably,markedly,marked,
risken	the risk,risk,
cliff	cliff,
nödvändigtvis	by necessity,necessarily,
knappast	hardly,dead,
inledning	introduction,
bysantinska	byzantine,
simpson	simpson,
tidning	newspaper,journal,
