vanligast	most	0	0	1	0
vanligast	most common	0	0	1	0
vanligast	most usual	0	0	1	0
nordisk	norse	0	0	1	0
nordisk	nordic	0	0	1	0
uppemot	almost	0	0	1	0
uppemot	up	0	0	1	0
förståelsen	the understanding	0	0	1	0
grundämnet	the element	0	0	1	0
grundämnet	element	0	0	1	0
stammarna	tribes	0	0	1	0
stammarna	strains	0	0	1	0
arternas	the species	0	0	1	0
arternas	species	0	0	1	0
uppleva	experience	0	0	1	1
jihad	johad	0	0	1	0
jihad	jihad	0	0	1	0
elva	eleven	0	0	1	1
invandrare	immigrants	0	0	1	0
invandrare	immigrant	0	0	1	1
luleå	luleå	0	0	1	0
albumet	album	0	0	1	0
besättningen	crew	0	0	1	0
albumen	the albums	0	0	1	0
albumen	albums	0	0	1	0
hermann	hermann	0	0	1	0
lord	lord	0	0	1	1
vann	won	0	0	1	0
lyckats	succeeded	0	0	1	0
dela	divide	0	0	1	1
dela	dividing	0	0	1	0
syrgas	oxygen	0	0	1	0
nuförtiden	nowadays	0	0	1	0
nuförtiden	today	0	0	1	0
regional	regional	0	0	1	1
upptar	occupies	0	0	1	0
portugals	portugals	0	0	1	0
portugals	portugal	0	0	1	0
dels	and	0	0	1	0
dels	both	0	0	1	0
dels	partly	0	0	1	1
skicklig	skillful	0	0	1	1
skicklig	proficient	0	0	1	1
skicklig	skilled; skillful	0	0	1	0
statlig	state	0	0	1	1
statlig	government	0	0	1	0
medelhavet	mediterranean sea	0	0	1	1
medelhavet	mediterranean	0	0	1	0
helsingborg	helsingborg	0	0	1	0
haber	haber	0	0	1	0
befogenheter	authorities	0	0	1	0
befogenheter	powers	0	0	1	0
triangelns	triangle	0	0	1	0
triangelns	the triangle's	0	0	1	0
kärnkraft	nuclear power	0	0	1	1
kärnkraft	nuclear	0	0	1	0
ögat	eye	0	0	1	0
urskilja	distinguish	0	0	1	1
urskilja	discern	0	0	1	1
sätter	place	0	0	1	0
sätter	puts	0	0	1	0
sätter	sets	0	0	1	0
sättet	manner	0	0	1	0
sättet	way	0	0	1	0
sättet	the way	0	0	1	0
sovjetisk	soviet	0	0	1	0
sovjetisk	sovjetic	0	0	1	0
sovjetisk	sovietic	0	0	1	0
miller	miller	0	0	1	0
hjärnans	the brain's	0	0	1	0
hjärnans	brain	0	0	1	0
sture	sture	0	0	1	0
målare	grinders	0	0	1	0
målare	painter	0	0	1	1
sammansatta	composite	0	0	1	0
sammansatta	composed	0	0	1	0
sammansatta	joined	0	0	1	0
grundämnen	elements	0	0	1	0
selassie	selassie	0	0	1	0
ungerns	hungary	0	0	1	0
ungerns	hungrarys	0	0	1	0
ungerns	hungary's	0	0	1	0
skilsmässa	divorce	0	0	1	1
hanar	males	0	0	1	0
makadam	congress	1	0	1	0
makadam	metal	1	0	1	1
makadam	macadam	1	1	0	1
makadam	tarmac	1	1	0	1
makadam	crushed rock	1	1	0	0
makadam	trip	1	0	1	0
breddgraden	latitude	0	0	1	0
breddgraden	parallel	0	0	1	0
fossil	fossil	0	0	1	1
punkt	item	0	0	1	1
punkt	point	0	0	1	1
filosofer	philosophers	0	0	1	0
filosofer	philosopher	0	0	1	0
aten	athens	0	0	1	0
biografi	biography	0	0	1	1
filosofen	the philosopher	0	0	1	0
regnskog	rain forest	0	0	1	0
regnskog	rainforest	0	0	1	1
herr	mister	0	0	1	1
herr	mr	0	0	1	0
misstänkta	suspected	0	0	1	0
misstänkta	suspect	0	0	1	0
kids	kids	0	0	1	0
demokratier	democracies	0	0	1	0
arabvärlden	the arab world	0	0	1	0
arabvärlden	arab world	0	0	1	0
naturen	the nature	0	0	1	0
naturen	nature	0	0	1	0
vicepresident	vice president	0	0	1	0
brottslighet	criminality	0	0	1	1
brottslighet	crime	0	0	1	1
miljarder	billion	0	0	1	0
miljarder	billions	0	0	1	0
karin	karin	0	0	1	0
systematiska	systematic	0	0	1	0
systematiska	systematical	0	0	1	0
unik	unique	0	0	1	1
norsk	norwegian	0	0	1	1
iis	ii's	0	0	1	0
marino	marino	0	0	1	0
västerländsk	western	0	0	1	1
hamas	hamas	0	0	1	0
större	greater	0	0	1	0
större	bigger	0	0	1	1
systematiskt	systematically	0	0	1	0
systematiskt	systematic	0	0	1	0
ansluta	join	0	0	1	0
ansluta	connect	0	0	1	1
närvarande	present (-ly)	0	0	1	0
närvarande	present	0	0	1	1
dna	dna	0	0	1	0
sjukdomen	disease	0	0	1	0
strikt	strict	0	0	1	0
hårdast	the most	0	0	1	0
hårdast	the hardest	0	0	1	0
hårdast	hardest	0	0	1	0
fuktiga	damp	0	0	1	0
fuktiga	futiga	0	0	1	0
fuktiga	damply	0	0	1	0
betraktats	considered	0	0	1	0
betraktats	been seen	0	0	1	0
betraktats	(been) viewed	0	0	1	0
music	music	0	0	1	0
dns	dns	0	0	1	0
fuktigt	moist	0	0	1	0
fuktigt	damp	0	0	1	0
fuktigt	humid	0	0	1	0
musik	music	0	0	1	1
mercurys	mercury's	0	0	1	0
mercurys	mercurys	0	0	1	0
bördiga	fertile	0	0	1	0
holm	holm	0	0	1	0
jordbävningar	earthquakes	0	0	1	0
politiker	politicians	0	0	1	0
politiker	politician	0	0	1	1
slutligen	back end	0	0	1	0
slutligen	at last	0	0	1	1
slutligen	finally	0	0	1	1
bulgariska	bulgarian	0	0	1	0
temperaturen	temperature	0	0	1	0
kalksten	limestone	0	0	1	1
särskilt	in particular	0	0	1	1
särskilt	particulary	0	0	1	0
särskilt	especially	0	0	1	1
högtider	holiday	0	0	1	0
högtider	feasts	0	0	1	0
teman	themes	0	0	1	0
teman	ternan	0	0	1	0
temperaturer	temperature	0	0	1	0
ofta	usually	0	0	1	0
ofta	often	0	0	1	1
särskild	specific	0	0	1	0
särskild	particular	0	0	1	1
avancerad	advanced	0	0	1	1
styrkan	strength; unit; force	0	0	1	0
styrkan	strength	0	0	1	0
väntade	expected	0	0	1	0
väntade	expected; were waiting	0	0	1	0
väntade	waited	0	0	1	0
befolkningsutveckling	population development	0	0	1	0
befolkningsutveckling	population growth	0	0	1	0
stommen	body	0	0	1	0
stommen	frame	0	0	1	0
stommen	the foundation	0	0	1	0
gjordes	made	0	0	1	0
gjordes	was	0	0	1	0
gjordes	was made	0	0	1	0
kapitalismen	capitalism	0	0	1	0
want	want	0	0	1	0
absoluta	absolute	0	0	1	0
korruptionsindex	corruption perceptions index	0	0	1	0
korruptionsindex	corruption index	0	0	1	0
domen	judgment	0	0	1	0
domen	verdict; judgement	0	0	1	0
näring	nutrition	0	0	1	1
hon	she	0	0	1	1
kallare	colder	0	0	1	0
hov	court	0	0	1	1
how	how	0	0	1	0
hot	hot	0	0	1	0
hos	with	0	0	1	1
hos	in; with	0	0	1	0
hos	of	0	0	1	0
folkmusik	folk music	0	0	1	1
könsorganen	sex organs	0	0	1	0
könsorganen	the reproductive organs	0	0	1	0
könsorganen	the genitals	0	0	1	0
koncentrationsläger	concentration	0	0	1	0
koncentrationsläger	concentration camp	0	0	1	1
koncentrationsläger	concentration camps; kz-camps	0	0	1	0
typen	model	0	0	1	0
typen	the type	0	0	1	0
typen	type	0	0	1	0
fylla	fill	0	0	1	1
inrikes	domestic	0	0	1	1
barbro	barbro	0	0	1	0
fyllt	filled	0	0	1	0
barney	barney	0	0	1	0
turkiet	turkey	0	0	1	1
turkiet	turklet	0	0	1	0
sankt	st.	0	0	1	1
sankt	sankt	0	0	1	0
typer	types	0	0	1	0
typer	characters	0	0	1	0
hisingen	hisingen	0	0	1	0
grekiska	greek	0	0	1	1
arbeten	works	0	0	1	0
deutsche	deutsche	0	0	1	0
köper	making	0	0	1	0
köper	buys	0	0	1	0
wind	wind	0	0	1	0
promemoria	short essay	1	0	1	0
promemoria		1	0	1	0
promemoria	memo	1	1	0	0
promemoria	memorandum	1	1	0	1
promemoria	aide-memoire	1	0	1	0
promemoria	stalin	1	0	1	0
promemoria	pm; memorandum	1	0	1	0
promemoria	pormemoria	1	0	1	0
promemoria	promemoria	1	0	1	0
vart	each	0	0	1	0
varv	revolutions	0	0	1	0
varv	dockyard	0	0	1	0
varv	shipbuilding	0	0	1	0
ormar	snakes	0	0	1	0
vars	whose	0	0	1	1
vars	who's	0	0	1	0
organismen	the organism	0	0	1	0
organismen	organism	0	0	1	0
vare	either	0	0	1	0
varg	wolf	0	0	1	1
organismer	organism	0	0	1	0
organismer	organisms	0	0	1	0
vara	be	0	0	1	1
omvandlas	convert	0	0	1	0
omvandlas	converted	0	0	1	0
mabel	mabel	0	0	1	0
belönades	rewarded	0	0	1	0
belönades	awarded	0	0	1	0
varm	hot	0	0	1	1
varm	warm	0	0	1	1
pojkvän	n/a	0	0	1	0
pojkvän	boyfriend	0	0	1	1
publicerade	published	0	0	1	0
klan	clan	0	0	1	1
okänd	unknown	0	0	1	1
vännen	the friend	0	0	1	0
vännen	friend	0	0	1	0
suveräna	terrific	0	0	1	0
suveräna	supreme	0	0	1	0
suveräna	sovereign	0	0	1	0
närmaste	nearest	0	0	1	0
närmaste	closest	0	0	1	0
nutida	present(-day); contemporary	0	0	1	0
nutida	present day	0	0	1	0
nutida	present	0	0	1	0
okänt	unknown	0	0	1	0
okänt	unkn	0	0	1	0
wales	wales	0	0	1	1
små	small	0	0	1	1
små	little	0	0	1	0
assyriska	assyrian	0	0	1	0
fil	master of	0	0	1	0
fil	file	0	0	1	1
hemlighet	secretly	0	0	1	0
hemlighet	darkness	0	0	1	1
suveränitet	sovereignty	0	0	1	1
euroområdet	eurozone	0	0	1	0
euroområdet	euro area	0	0	1	0
euroområdet	convergence report	0	0	1	0
silver	silver	0	0	1	1
utvecklat	developed	0	0	1	0
utvecklat	evolved	0	0	1	0
tyder	indicates	0	0	1	0
utvecklar	develops	0	0	1	0
utvecklar	development speaker	0	0	1	0
utvecklas	development	0	0	1	0
terrorister	terrorists	0	0	1	0
tingslag	leet	0	0	1	0
tingslag	things type	0	0	1	0
debut	debut	0	0	1	1
utveckling	development	0	0	1	1
utvecklad	developed	0	0	1	0
påven	the pope	0	0	1	0
påven	paven	0	0	1	0
påven	pope	0	0	1	0
köpenhamn	copenhagen	0	0	1	1
ingrid	ingrid	0	0	1	0
därefter	then	0	0	1	1
därefter	thereafter	0	0	1	1
likväl	nevertheless	0	0	1	1
likväl	still	0	0	1	0
likväl	as well	0	0	1	0
talade	spoken	0	0	1	0
talade	spoke	0	0	1	0
sapiens	sapiens	0	0	1	0
angola	angola	0	0	1	1
treenighetsläran	doctrine of the holy trinity	0	0	1	0
treenighetsläran	trinity	0	0	1	0
treenighetsläran	school of trinity	0	0	1	0
serier	comics	0	0	1	0
serier	series	0	0	1	0
allan	allan	0	0	1	0
utvecklandet	development	0	0	1	0
serien	series	0	0	1	0
serien	the series	0	0	1	0
arab	arab	0	0	1	1
truman	truman	0	0	1	0
uppmärksammades	attention	0	0	1	0
uppmärksammades	drew attention	0	0	1	0
varken	neither	0	0	1	1
varken	either	0	0	1	0
kontrollerade	controlled	0	0	1	1
slovenien	slovenia	0	0	1	1
slovenien	slovenian	0	0	1	0
innehållande	containing	0	0	1	1
innehållande	including	0	0	1	0
foundation	foundation	0	0	1	0
snarare	rather	0	0	1	1
nuvarande	current	0	0	1	1
anarkister	anarchists	0	0	1	0
metallica	metallica	0	0	1	0
arbetsplats	work	0	0	1	0
arbetsplats	workplace	0	0	1	0
sannolikt	probably	0	0	1	0
sannolikt	probable	0	0	1	0
att	to	0	0	1	1
att	that	0	0	1	1
atp	atp	0	0	1	0
sydost	south east	0	0	1	0
sydost	southeast	0	0	1	0
landområden	land	0	0	1	0
landområden	land areas	0	0	1	0
givetvis	course	0	0	1	0
givetvis	naturally	0	0	1	1
debatten	debate	0	0	1	0
debatten	the debate	0	0	1	0
affärer	business	0	0	1	0
tecknade	cartoon (-s)	0	0	1	0
tecknade	cartoon	0	0	1	0
tecknade	drew	0	0	1	0
service	service	0	0	1	1
xii	xii	0	0	1	0
xis	the eleventh's	0	0	1	0
master	masters	0	0	1	0
master	master	0	0	1	0
bitter	bitter	0	0	1	1
senaten	senate	0	0	1	0
senaten	the senate	0	0	1	0
undantaget	except	0	0	1	0
begärde	called	0	0	1	0
begärde	demanded	0	0	1	0
placerade	put	0	0	1	0
placerade	placed	0	0	1	0
placerade	placed (in)	0	0	1	0
nirvana	nirvana	0	0	1	1
susan	susan	0	0	1	0
ahmed	ahmed	0	0	1	0
skatter	taxes	0	0	1	0
upphov	origin	0	0	1	1
upphov	source	0	0	1	1
upphov	rise	0	0	1	0
tyckte	thought	0	0	1	0
tyckte	found	0	0	1	0
tyckte	find	0	0	1	0
tree	tree	0	0	1	0
gator	streets	0	0	1	0
nations	nations	0	0	1	0
nations	nation	0	0	1	0
trey	trey	0	0	1	0
varje	each	0	0	1	1
utformningen	the layout	0	0	1	0
utformningen	layout	0	0	1	0
utformningen	the design	0	0	1	0
östtyska	east german	0	0	1	0
tretton	thirteen	0	0	1	1
obligatorisk	obligatory	0	0	1	1
obligatorisk	mandatory	0	0	1	1
järnväg	railroad	0	0	1	1
järnväg	rail	0	0	1	1
järnväg	railway	0	0	1	1
assistent	assistant	0	0	1	1
kriterierna	criteria	0	0	1	0
boston	boston	0	0	1	1
dricker	drinking	0	0	1	0
dricker	drink	0	0	1	0
dricker	drinks	0	0	1	0
filosofisk	philosophical	0	0	1	0
filosofisk	philosophic	0	0	1	1
sågs	observed	0	0	1	0
sågs	seen	0	0	1	0
sågs	was observed	0	0	1	0
halva	half	0	0	1	1
joakim	joakim	0	0	1	0
trakten	the region	0	0	1	0
trakten	region	0	0	1	0
trakten	area	0	0	1	0
fasta	solid	0	0	1	0
fasta	firm; set; solid; fast; fasting	0	0	1	0
kroatien	croatia	0	0	1	1
händerna	the hands	0	0	1	0
händerna	hands	0	0	1	0
konstnärlig	art	0	0	1	0
konstnärlig	artistic	0	0	1	1
krigsmakt	military power	0	0	1	0
krigsmakt	armed forces	0	0	1	0
fastän	although	0	0	1	1
skaffa	obtain	0	0	1	1
skaffa	gain	0	0	1	0
skaffa	get	0	0	1	1
spelningar	tour	0	0	1	0
spelningar	gigs	0	0	1	0
öar	islets	0	0	1	0
öar	islands	0	0	1	0
himlen	heaven	0	0	1	0
himlen	although the sky	0	0	1	0
utgåva	edition	0	0	1	1
utgåva	issue	0	0	1	1
bedrivs	conducted	0	0	1	0
katalonien	catalonia	0	0	1	0
konserthus	concert hall	0	0	1	0
konserthus	concert	0	0	1	0
victoria	victoria	0	0	1	0
gallagher	gallagher	0	0	1	0
medlemsstaterna	member	0	0	1	0
medlemsstaterna	member states	0	0	1	0
anteckningar	notes	0	0	1	0
bedriva	carry	0	0	1	0
bedriva	prosecute	0	0	1	1
eftersom	while	0	0	1	0
eftersom	because	0	0	1	0
thriller	thriller	0	0	1	1
annars	else	0	0	1	1
singer	singer	0	0	1	0
morgon	tomorrow	0	0	1	0
morgon	morning	0	0	1	1
förväxla	confuse	0	0	1	1
förväxla	mistake	0	0	1	0
arkitektur	architecture	0	0	1	1
professor	professor	0	0	1	1
camp	camp	0	0	1	0
nederbörden	precipitation	0	0	1	0
nederbörden	the precipitation	0	0	1	0
mängd	volume	0	0	1	0
mängd	amount	0	0	1	1
mängd	laden	0	0	1	0
grovt	heavy	0	0	1	0
grovt	rough	0	0	1	0
grovt	roughly	0	0	1	0
passerade	passed	0	0	1	0
singel	single	0	0	1	0
inspelning	recording	0	0	1	1
ungar	kids	0	0	1	0
ungar	babies	0	0	1	0
ungar	kids; offsprings; young	0	0	1	0
bomb	bomb	0	0	1	1
bandmedlemmar	band members	0	0	1	0
nacka	nacka	0	0	1	0
pris	price	0	0	1	1
pris	prize	0	0	1	1
teater	theatre; theater	0	0	1	0
teater	theater	0	0	1	1
louise	louis	0	0	1	0
louise	louise	0	0	1	0
lönneberga	lönneberga	0	0	1	0
lönneberga	lonneberga	0	0	1	0
buss	bus	0	0	1	1
delats	divided	0	0	1	0
delats	been awarded	0	0	1	0
rico	rico	0	0	1	0
bush	bush	0	0	1	0
rice	rice	0	0	1	0
mottog	received	0	0	1	0
lastbilar	truck	0	0	1	0
lastbilar	trucks	0	0	1	0
storbritanniens	united kingdom	0	0	1	0
storbritanniens	uk	0	0	1	0
ämnena	subjects	0	0	1	0
ämnena	the elements	0	0	1	0
ämnena	substances	0	0	1	0
kompositör	composer	0	0	1	1
digerdöden	black death	0	0	1	0
digerdöden	digerdoden	0	0	1	0
digerdöden	the black death	0	0	1	0
metoder	methods	0	0	1	0
platt	flat	0	0	1	1
platt	plate	0	0	1	0
metoden	the method	0	0	1	0
dansk	danish	0	0	1	1
plats	spot	0	0	1	0
plats	place	0	0	1	1
plats	place; position	0	0	1	0
bensin	gasoline	0	0	1	1
lyssna	listening	0	0	1	0
lyssna	listen	0	0	1	1
begravning	funeral	0	0	1	1
stödde	supported	0	0	1	0
medfört	resulted	0	0	1	0
medfört	led to	0	0	1	0
hantverk	crafting	0	0	1	0
hantverk	crafts	0	0	1	1
kallt	cold	0	0	1	0
kallt	coldly	0	0	1	1
dröja	take	0	0	1	0
dröja	wait	0	0	1	1
framfört	expressed	0	0	1	0
framfört	presented	0	0	1	0
uppgift	task	0	0	1	1
uppgift	data	0	0	1	0
övergår	surpasses	0	0	1	0
övergår	released	0	0	1	0
övergår	exceed	0	0	1	0
framförs	is presented	0	0	1	0
framförs	performed	0	0	1	0
kalle	kalle	0	0	1	0
höst	autumn	0	0	1	1
höst	fall	0	0	1	1
kalla	cold	0	0	1	0
ovtjarka	ovtjarka	0	0	1	0
ovtjarka	caucasian shepherd dog	0	0	1	0
händelsehorisonten	event horizon	0	0	1	0
händelsehorisonten	the event horizon	0	0	1	0
händelsehorisonten	place else horizon	0	0	1	0
blev	became	0	0	1	0
blev	was	0	0	1	0
etik	ethics	0	0	1	1
flagga	flag	0	0	1	1
skulle	could	0	0	1	0
skulle	would	0	0	1	1
skriva	write	0	0	1	1
bygger	based	0	0	1	0
bygger	(is) building (on)	0	0	1	0
erövrade	conquered	0	0	1	0
arlanda	arlanda	0	0	1	0
skrivs	written	0	0	1	0
skrivs	printed	0	0	1	0
våningar	floors	0	0	1	0
våningar	storeys	0	0	1	0
hedersdoktor	honorary doctor	0	0	1	1
hedersdoktor	honorary degree	0	0	1	0
hedersdoktor	honorary doctorate	0	0	1	0
manson	manson	0	0	1	0
dröjde	slow	0	0	1	0
dröjde	was not until	0	0	1	0
dröjde	not until	0	0	1	0
wikipedia	wikipedia	0	0	1	0
sundsvalls	sundsvall	0	0	1	0
sundsvalls	(city of) sundsvall's	0	0	1	0
ägna	devote	0	0	1	1
ägna	spend	0	0	1	0
ägna	baiting	0	0	1	0
figur	figure	0	0	1	1
sista	last	0	0	1	1
siste	lattermost	0	0	1	1
siste	last	0	0	1	0
pirate	pirate	0	0	1	0
ringa	call	0	0	1	1
rollen	role	0	0	1	0
rollen	the role	0	0	1	0
henrik	henrik	0	0	1	0
tropisk	tropical	0	0	1	1
lanserades	launched	0	0	1	0
lanserades	was launched	0	0	1	0
bestämma	determining	0	0	1	0
bestämma	decide	0	0	1	1
tilldelades	awarded	0	0	1	0
kommunikation	communication	0	0	1	1
kommunikation	communications	0	0	1	0
roller	roles	0	0	1	0
kloster	monastery	0	0	1	1
huvudet	head	0	0	1	0
huvudet	the head	0	0	1	0
krönika	chronicle	0	0	1	1
country	country	0	0	1	0
gärningsmannen	perpetrator; offender	0	0	1	0
gärningsmannen	the offender	0	0	1	0
gärningsmannen	culprit	0	0	1	0
pitt	pitt	0	0	1	0
edgar	edgar	0	0	1	0
nordiska	nordic	0	0	1	1
rädda	save	0	0	1	1
rädda	lot of	0	0	1	0
förstnämnda	first-named	0	0	1	0
förstnämnda	aforementioned	0	0	1	0
förstnämnda	first named	0	0	1	0
besserwisser	a	1	0	1	0
besserwisser	pundit	1	0	1	0
besserwisser	give	1	0	1	0
besserwisser	between	1	0	1	0
besserwisser	exact: better knower; equivalent: know-it-all	1	0	1	0
besserwisser	know it all	1	1	0	0
besserwisser	smartass	1	0	1	0
besserwisser	know-all	1	1	0	1
besserwisser	know-it-all	1	1	0	0
besserwisser	bewiseacre	1	0	1	0
besserwisser	besserwisser	1	1	0	0
besserwisser	wiseacre	1	1	0	1
anordnas	provided	0	0	1	0
anordnas	arranged	0	0	1	0
anordnas	organised	0	0	1	0
nordiskt	nordic	0	0	1	0
genus	gender	0	0	1	1
genus	genus	0	0	1	0
logik	logic	0	0	1	1
summan	sum	0	0	1	0
summan	the sum	0	0	1	0
igelkotten	the hedgehog	0	0	1	0
igelkotten	hedgehog	0	0	1	0
förgäves	in vain	0	0	1	1
folkmordet	genocide	0	0	1	0
färre	fewer	0	0	1	1
färre	less	0	0	1	0
rumänien	romania	0	0	1	0
brännvin	schnaps	0	0	1	0
brännvin	aquavit	0	0	1	0
äktenskapet	marriage	0	0	1	0
uttal	pronunciation	0	0	1	1
uttal	pronounciation	0	0	1	0
analytisk	analytical	0	0	1	1
afrikanska	afrikanska	0	0	1	0
afrikanska	african	0	0	1	0
fra	fra	0	0	1	0
union	union	0	0	1	1
fri	free	0	0	1	1
tiotusentals	tens of thousands	0	0	1	0
operationer	operations	0	0	1	1
socialistiskt	socialistic	0	0	1	0
socialistiskt	socialist	0	0	1	0
fru	madam	0	0	1	0
fru	mrs.	0	0	1	1
fru	wife	0	0	1	1
verktyg	tool	0	0	1	1
verktyg	tools	0	0	1	0
socialistiska	socialistic	0	0	1	0
socialistiska	socialist	0	0	1	0
life	life	0	0	1	0
snittet	average	0	0	1	0
snittet	the intersection	0	0	1	0
snittet	the average	0	0	1	0
arkiv	archives	0	0	1	1
arkiv	archive	0	0	1	0
dave	dave	0	0	1	0
kometer	comets	0	0	1	0
chile	chile	0	0	1	1
motorvägen	motorway	0	0	1	0
motorvägen	highway	0	0	1	0
chili	chili	0	0	1	1
hålls	is held	0	0	1	0
hålls	maintaned	0	0	1	0
hålls	maintained	0	0	1	0
intag	intake	0	0	1	1
slutliga	evenutal	0	0	1	0
slutliga	final	0	0	1	0
slutliga	ultimate	0	0	1	0
frankrikes	france's	0	0	1	0
frankrikes	frances	0	0	1	0
önskemål	desire	0	0	1	1
önskemål	requests	0	0	1	0
önskemål	demands	0	0	1	0
castro	castro	0	0	1	0
hålla	hold	0	0	1	1
hålla	keep	0	0	1	1
klarade	made it	0	0	1	0
klarade	passed	0	0	1	0
organisera	organize	0	0	1	1
organisera	organizing	0	0	1	0
kontraktet	the contract	0	0	1	0
kontraktet	contract	0	0	1	0
tintin	tintin	0	0	1	0
k	k	0	0	1	0
erövra	conquer	0	0	1	1
fyllde	completed	0	0	1	0
fyllde	filled	0	0	1	0
brister	failures	0	0	1	0
brister	inabilities	0	0	1	0
desto	the	0	0	1	0
desto	ever	0	0	1	0
kurderna	kurdish	0	0	1	0
kurderna	kurds	0	0	1	0
player	player	0	0	1	0
fascismen	the fascism	0	0	1	0
fascismen	fascism	0	0	1	0
bristen	lack of	0	0	1	0
bristen	lack	0	0	1	0
folkmängd	population size	0	0	1	0
folkmängd	population	0	0	1	1
madonna	madonna	0	0	1	1
räckte	enough	0	0	1	0
räckte	handed	0	0	1	1
azidgrupp	azido group	1	0	1	0
azidgrupp	azide	1	1	0	0
azidgrupp	lost	1	0	1	0
azidgrupp	amide	1	0	1	0
azidgrupp	azite group	1	0	1	0
azidgrupp	azid group	1	1	0	0
azidgrupp	azide group	1	1	0	0
azidgrupp	azidgrupp	1	0	1	0
memorial	memorial	0	0	1	0
serbisk	serbian	0	0	1	1
vrida	twist	0	0	1	1
vrida	turn	0	0	1	1
vrida	turning	0	0	1	0
foton	images	0	0	1	0
foton	photos	0	0	1	0
omkring	surrounding	0	0	1	0
omkring	about	0	0	1	1
omkring	around	0	0	1	1
agnetha	agnetha	0	0	1	0
european	european	0	0	1	0
än	than	0	0	1	1
än	yet	0	0	1	1
materiell	materiell	0	0	1	0
materiell	material	0	0	1	1
funktionen	function	0	0	1	0
funktionen	the function	0	0	1	0
josef	joseph	0	0	1	0
josef	josef	0	0	1	0
topp	top	0	0	1	1
linné	linen	0	0	1	0
linné	linneus	0	0	1	0
linné	temperature	0	0	1	0
tunn	thin	0	0	1	1
funktioner	functions	0	0	1	0
funktioner	features	0	0	1	0
synder	sins	0	0	1	0
tung	heavy	0	0	1	1
obligatoriskt	obligatory	0	0	1	0
obligatoriskt	mandatory	0	0	1	0
efterföljare	following	0	0	1	0
efterföljare	follower	0	0	1	1
efterföljare	successors	0	0	1	0
finska	finnish	0	0	1	0
lucas	lucas	0	0	1	0
kampanj	campaign	0	0	1	1
centraleuropa	central europe	0	0	1	0
ansågs	was	0	0	1	0
ansågs	seemed	0	0	1	0
gudinnan	goddess	0	0	1	0
gudinnan	the godess	0	0	1	0
grundlag	constitution	0	0	1	1
misslyckade	failed	0	0	1	0
manteln	the mantle	0	0	1	0
manteln	mantle	0	0	1	0
koloniseringen	the colonization	0	0	1	0
koloniseringen	colonization	0	0	1	0
fortplantning	reproduction	0	0	1	1
fortplantning	sex	0	0	1	0
grönsaker	vegetables	0	0	1	1
krigsmakten	war food	0	0	1	0
krigsmakten	armed forces	0	0	1	0
birmingham	birmingham	0	0	1	1
lasse	lasse	0	0	1	0
kommunal	communal	0	0	1	1
kommunal	municipal	0	0	1	1
givit	gave	0	0	1	0
matteus	matthew	0	0	1	0
matteus	matteus	0	0	1	0
han	he	0	0	1	1
grafit	graphite	0	0	1	1
bnp	gdp	0	0	1	0
bnp	gnp	0	0	1	0
fysikaliska	physical	0	0	1	0
muhammeds	mohammed's	0	0	1	0
muhammeds	muhammad	0	0	1	0
muhammeds	muhammed's	0	0	1	0
huvud	head	0	0	1	1
huvud	main	0	0	1	0
hette	name was	0	0	1	0
hette	hatte	0	0	1	0
hette	named	0	0	1	0
lunginflammation	pneumonia	0	0	1	1
har	is	0	0	1	0
har	has	0	0	1	0
har	have	0	0	1	0
hat	hatred	0	0	1	1
hav	seas	0	0	1	0
hav	sea	0	0	1	1
hav	ocean	0	0	1	1
kön	gender	0	0	1	1
kön	sex	0	0	1	1
underliggande	underlying	0	0	1	1
svensson	svensson	0	0	1	0
svensson	smith	0	0	1	0
narkotika	drug	0	0	1	1
narkotika	narcotics	0	0	1	0
livsstil	life style	0	0	1	0
livsstil	lifestyle	0	0	1	0
älskar	loves	0	0	1	0
kör	run	0	0	1	0
melodifestivalen	eurovision song contest	0	0	1	0
melodifestivalen	music festival	0	0	1	0
köp	purchase	0	0	1	1
county	county	0	0	1	0
bobby	bobby	0	0	1	0
tågen	train	0	0	1	0
tågen	the trains	0	0	1	0
sedlar	bills	0	0	1	0
alice	alice	0	0	1	0
kust	coastal	0	0	1	0
kust	coast	0	0	1	1
residensstad	city of residence	0	0	1	0
residensstad	county seat	0	0	1	0
tåget	train	0	0	1	0
tåget	the train	0	0	1	0
moral	morality	0	0	1	1
sebastian	sebastian	0	0	1	0
grannländer	neighbors	0	0	1	0
grannländer	neighboring countries	0	0	1	0
grannländer	neighboring lander	0	0	1	0
ola	ola	0	0	1	0
old	old	0	0	1	0
interstellära	interstellar	0	0	1	0
people	people	0	0	1	0
billboard	billboard	0	0	1	0
parlamentarisk	parliamentary	0	0	1	0
delade	shared	0	0	1	0
delade	divided	0	0	1	0
delade	split	0	0	1	0
rörelserna	the movements	0	0	1	0
rörelserna	movement	0	0	1	0
kulmen	culmination	0	0	1	1
kulmen	the acme	0	0	1	0
kulmen	peak	0	0	1	0
fot	foot	0	0	1	1
fot	ft	0	0	1	0
föga	little	0	0	1	1
föga	hardly; little	0	0	1	0
for	for	0	0	1	0
varierande	variable	0	0	1	1
varierande	varied	0	0	1	1
varierande	varying	0	0	1	1
fox	fox	0	0	1	0
utser	chooses	0	0	1	0
utser	appoints	0	0	1	0
utses	is appointed	0	0	1	0
utses	designated	0	0	1	0
utses	appointed	0	0	1	0
akademi	academy	0	0	1	1
framstående	prominent	0	0	1	0
bokstäverna	the letters	0	0	1	0
bokstäverna	letters	0	0	1	0
järnvägsnätet	railroad network	0	0	1	0
järnvägsnätet	rail	0	0	1	0
myndigheter	authorities	0	0	1	0
myndigheter	agencies	0	0	1	0
annan	another	0	0	1	0
inkomstkälla	income cold	0	0	1	0
inkomstkälla	was added to cold	0	0	1	0
inkomstkälla	source of income	0	0	1	1
neptunus	neptunes	0	0	1	0
neptunus	neptune	0	0	1	1
stefan	stefan	0	0	1	0
översättningen	translation	0	0	1	0
översättningen	the translation	0	0	1	0
binder	bind	0	0	1	0
binder	tie	0	0	1	0
olympiska	olympic	0	0	1	0
älg	elk	0	0	1	1
älg	moose	0	0	1	1
myndigheten	the authority	0	0	1	0
myndigheten	authority	0	0	1	0
annat	alia	0	0	1	0
annat	other	0	0	1	1
annat	other; another	0	0	1	0
beräkna	calculated	0	0	1	0
beräkna	calculate	0	0	1	1
army	army	0	0	1	0
o	oh	0	0	1	0
mynnar	opening	0	0	1	0
klubben	club	0	0	1	0
nixon	nixon	0	0	1	0
tillverkare	producer	0	0	1	0
tillverkare	manufacturer	0	0	1	1
delvis	partly	0	0	1	1
delvis	partial	0	0	1	1
delvis	partially	0	0	1	1
psykiska	psychic	0	0	1	0
psykiska	mental	0	0	1	0
material	material	0	0	1	1
material	materials	0	0	1	0
marshall	marshall	0	0	1	0
som	as	0	0	1	1
som	which	0	0	1	1
sol	sun	0	0	1	1
lagliga	legal	0	0	1	0
lagliga	lawful	0	0	1	0
son	son	0	0	1	1
psykiskt	psychic	0	0	1	0
psykiskt	mentally	0	0	1	0
västindien	caribbean	0	0	1	0
västindien	west india	0	0	1	0
skådespelarna	actors	0	0	1	0
skådespelarna	period players	0	0	1	0
fci	fci	0	0	1	0
ingående	input	0	0	1	0
ingående	in depth	0	0	1	0
ingående	enter into	0	0	1	0
delarna	the parts	0	0	1	0
delarna	parts	0	0	1	0
alltså	so	0	0	1	1
alltså	therefore	0	0	1	0
alltså	really	0	0	1	0
artikeln	the article	0	0	1	0
hantera	handle	0	0	1	1
nova	nova	0	0	1	0
joseph	joseph	0	0	1	0
böhmen	bohemia	0	0	1	1
jane	jane	0	0	1	0
happy	happy	0	0	1	0
offer	victims	0	0	1	1
offer	victim	0	0	1	1
verde	verde	0	0	1	0
enighet	unity	0	0	1	1
drabbat	affected	0	0	1	0
gymnasiet	high school	0	0	1	0
gymnasiet	gymnasium	0	0	1	0
drabbar	affect	0	0	1	0
drabbar	troubles	0	0	1	0
drabbar	afflict	0	0	1	0
polska	polish	0	0	1	1
mörkt	dark	0	0	1	0
syften	purpose	0	0	1	0
pest	plague	0	0	1	1
syftet	purpose	0	0	1	0
tänderna	tandem	0	0	1	0
tänderna	teeh	0	0	1	0
tänderna	teeth	0	0	1	0
mörka	dark	0	0	1	0
mörka	morka	0	0	1	0
fansen	fans	0	0	1	0
fansen	the fan	0	0	1	0
moderna	modern	0	0	1	0
liberal	liberal	0	0	1	1
konung	king	0	0	1	1
lunds	lund's	0	0	1	0
lunds	lund	0	0	1	0
modernt	modern	0	0	1	0
länder	states	0	0	1	0
länder	countries	0	0	1	0
ericsson	ericsson	0	0	1	0
nämnts	mentioned	0	0	1	0
nämnts	above	0	0	1	0
nordväst	north west	0	0	1	0
nordväst	northwest	0	0	1	0
elektromagnetisk	electromagnetic	0	0	1	0
huvudperson	main person; main character	0	0	1	0
huvudperson	protagonist	0	0	1	1
huvudperson	main character	0	0	1	0
oväntat	unexpectedly	0	0	1	1
oväntat	unexpected	0	0	1	0
dotter	daughter	0	0	1	1
protester	protests	0	0	1	0
republik	republic	0	0	1	1
roll	role	0	0	1	1
olja	oil	0	0	1	1
föreslår	proposes	0	0	1	0
föreslår	suggests	0	0	1	0
föreslår	suggest	0	0	1	0
reggae	reggae	0	0	1	0
avskaffades	was abolished	0	0	1	0
avskaffades	abolished	0	0	1	0
runda	round	0	0	1	1
palme	palme	0	0	1	0
vintrarna	the winters	0	0	1	0
vintrarna	winters	0	0	1	0
modell	model	0	0	1	1
rolling	rolling	0	0	1	0
utbildade	formed	0	0	1	0
utbildade	educated	0	0	1	0
danske	danish	0	0	1	0
danske	dane	0	0	1	0
aragorn	aragorn	0	0	1	0
avståndet	distance	0	0	1	0
avståndet	the distance	0	0	1	0
danska	danish	0	0	1	1
motståndaren	adversary	0	0	1	0
motståndaren	the opponent	0	0	1	0
motståndaren	opponent	0	0	1	0
povel	povel	0	0	1	0
laddade	charged	0	0	1	0
perioden	period	0	0	1	0
perioden	time	0	0	1	0
trettio	thirty	0	0	1	1
perioder	periods; episodes	0	0	1	0
perioder	period	0	0	1	0
perioder	periods	0	0	1	0
time	time	0	0	1	0
östergötland	Östergötland	0	0	1	0
östergötland	east gothland	0	0	1	0
skatt	tax	0	0	1	1
sträckte	extended	0	0	1	0
oss	center	0	0	1	0
oss	us	0	0	1	1
ost	cheese	0	0	1	1
uppgifter	information	0	0	1	1
uppgifter	tasks	0	0	1	0
uppgifter	data	0	0	1	0
avalanche	avalanche	0	0	1	0
uppgiften	the task	0	0	1	0
uppgiften	task	0	0	1	0
atombomben	atom bomb	0	0	1	0
atombomben	atomic bomb	0	0	1	0
atombomben	the nuclear bomb	0	0	1	0
traditionell	traditional	0	0	1	1
traditionell	conventional	0	0	1	0
efterfrågan	the demand	0	0	1	0
efterfrågan	demand	0	0	1	1
inkomst	income	0	0	1	1
machu	machu	0	0	1	0
vet	know	0	0	1	0
öga	eye	0	0	1	1
hjälpmedel	aid	0	0	1	1
hjälpmedel	means agent	0	0	1	0
hjälpmedel	resources	0	0	1	0
intresserade	interested	0	0	1	0
regissören	director	0	0	1	0
vem	who	0	0	1	1
åtta	eight	0	0	1	1
bosnien	bosnian	0	0	1	0
bosnien	bosnia	0	0	1	1
musikstilar	music genres	0	0	1	0
musikstilar	music	0	0	1	0
individer	individuals	0	0	1	0
individer	subjects	0	0	1	0
choice	choice	0	0	1	0
individen	the individual	0	0	1	0
individen	individual	0	0	1	0
skillnaderna	the differences	0	0	1	0
skillnaderna	differences	0	0	1	0
kusterna	the coasts	0	0	1	0
kusterna	coasts	0	0	1	0
initiativ	initiative	0	0	1	1
däggdjur	mammalian	0	0	1	0
däggdjur	mammal	0	0	1	1
hörde	heard	0	0	1	0
inhemska	native	0	0	1	0
smålands	smaland's	0	0	1	0
smålands	småland	0	0	1	0
energin	the energy	0	0	1	0
energin	energy	0	0	1	0
oppositionen	opposition	0	0	1	0
modersmål	native language	0	0	1	1
modersmål	mother tongue	0	0	1	1
team	team	0	0	1	1
uppskattningsvis	estimated	0	0	1	0
uppskattningsvis	approximately	0	0	1	0
uppskattningsvis	an estimated	0	0	1	0
be	be	0	0	1	0
fängelse	prison	0	0	1	1
scen	scene	0	0	1	1
scen	stage	0	0	1	1
tros	belived	0	0	1	0
tros	believed	0	0	1	0
firandet	the celebration	0	0	1	0
firandet	celebrate	0	0	1	0
låtar	songs	0	0	1	0
målen	cases	0	0	1	0
målen	goals	0	0	1	0
elton	elton	0	0	1	0
elton	tone	0	0	1	0
kunskapen	the knowledge	0	0	1	0
kunskapen	knowledge	0	0	1	0
strävar	striving; aiming (to; for)	0	0	1	0
strävar	strives	0	0	1	0
beskydd	conservation	0	0	1	0
beskydd	protection	0	0	1	1
axel	axel	0	0	1	0
strävan	will	0	0	1	0
strävan	the quest	0	0	1	0
strävan	endeavor	0	0	1	1
bosatte	settled	0	0	1	0
kunskaper	knowledge	0	0	1	1
bosatta	residents	0	0	1	0
bosatta	settled	0	0	1	0
västeuropeiska	western european	0	0	1	0
västeuropeiska	living	0	0	1	0
kusten	the coast	0	0	1	0
kusten	coast	0	0	1	0
katter	cats	0	0	1	0
katter	cat	0	0	1	0
provinserna	provinces	0	0	1	0
provinserna	the provinces	0	0	1	0
galileo	galileo	0	0	1	0
vintertid	winter-time	0	0	1	0
vintertid	winter	0	0	1	0
budskapet	the  message	0	0	1	0
budskapet	the message	0	0	1	0
budskapet	message	0	0	1	0
katten	the cat	0	0	1	0
katten	cat	0	0	1	0
huvudsakliga	main	0	0	1	0
studien	study	0	0	1	0
studien	the study	0	0	1	0
använder	using	0	0	1	0
använder	uses	0	0	1	0
användes	was used	0	0	1	0
användes	used	0	0	1	0
överallt	in all	0	0	1	0
överallt	everywhere	0	0	1	1
överallt	overall; everywhere	0	0	1	0
landslag	national team	0	0	1	0
studiet	study	0	0	1	0
studiet	the study	0	0	1	0
studier	studies	0	0	1	0
resande	travelers	0	0	1	0
resande	travelling	0	0	1	1
love	love	0	0	1	0
beläget	located	0	0	1	0
beläget	base	0	0	1	0
tidskriften	the magazine	0	0	1	0
tidskriften	magazine	0	0	1	0
kommit	to be	0	0	1	0
kommit	come	0	0	1	0
rocksångare	rock singers	0	0	1	0
rocksångare	rock singer	0	0	1	0
presenterade	travel related	0	0	1	0
presenterade	presented	0	0	1	0
canis	canis	0	0	1	0
sprids	spreading	0	0	1	0
sprids	spreads	0	0	1	0
samlat	collected	0	0	1	0
samlat	single	0	0	1	0
samlat	gathered	0	0	1	0
samlar	collect	0	0	1	0
samlar	salmar	0	0	1	0
samlar	collectors	0	0	1	0
positiva	positive	0	0	1	0
vuxna	adult	0	0	1	0
emellan	a	0	0	1	0
emellan	inbetween; between	0	0	1	0
emellan	between	0	0	1	1
neologi	neologism	1	0	1	0
neologi		1	0	1	0
neologi	neology	1	1	0	0
neologi	plans	1	0	1	0
neologi	projected	1	0	1	0
neologi	neologi	1	0	1	0
neologi	planned	1	0	1	0
neologi	a new logical	1	1	0	0
neologi	girl	1	0	1	0
judarna	the jews	0	0	1	0
judarna	jews	0	0	1	0
judarna	therefore	0	0	1	0
positivt	positive	0	0	1	0
samlag	intercourse	0	0	1	0
stärktes	was strengthened	0	0	1	0
stärktes	strengthened	0	0	1	0
stärktes	was strenghten	0	0	1	0
ökade	increased	0	0	1	0
påståenden	claims	0	0	1	0
påståenden	assertions	0	0	1	0
kött	meat	0	0	1	1
kött	cones	0	0	1	0
dagars	day's	0	0	1	0
dagars	day	0	0	1	0
dagars	days	0	0	1	0
relationerna	the relationships	0	0	1	0
relationerna	relations	0	0	1	0
stjärnorna	stars	0	0	1	0
stjärnorna	the stars	0	0	1	0
tabellen	table	0	0	1	0
tabellen	the chart	0	0	1	0
tabellen	table; list	0	0	1	0
soldaterna	soldiers	0	0	1	0
soldaterna	the soldiers	0	0	1	0
straffet	penalty	0	0	1	0
straffet	the punishment	0	0	1	0
kunskap	knowledge	0	0	1	1
sönder	broken	0	0	1	1
sönder	probes	0	0	1	0
phoebe	phoebe	0	0	1	0
phoebe	hoebe	0	0	1	0
förde	forde	0	0	1	0
förde	led	0	0	1	0
förde	out	0	0	1	0
stigande	rising	0	0	1	1
stigande	up	0	0	1	0
så	as	0	0	1	1
så	so	0	0	1	1
locka	attract	0	0	1	0
locka	tempt	0	0	1	1
gäller	of	0	0	1	0
gäller	refer to	0	0	1	0
gäller	grating	0	0	1	0
locke	locke	0	0	1	0
inkluderade	included	0	0	1	0
sångare	singer	0	0	1	1
kretsar	circuits	0	0	1	0
kretsar	circles	0	0	1	0
kretsar	circuitry	0	0	1	0
väsentligt	substantially	0	0	1	0
väsentligt	relevant	0	0	1	0
utnyttjade	utilized	0	0	1	0
utnyttjade	used	0	0	1	0
svenskar	swedish	0	0	1	0
svenskar	swedes	0	0	1	0
milda	mild	0	0	1	0
skikt	layers	0	0	1	0
skikt	layer	0	0	1	1
svenskan	swedish	0	0	1	0
svenskan	the swede	0	0	1	0
storleken	size	0	0	1	0
trigonometriska	trigonometric	0	0	1	0
levande	live	0	0	1	1
riksdagen	parliament	0	0	1	0
riksdagen	the parliament	0	0	1	0
gigantiska	gigantic	0	0	1	0
gigantiska	giant	0	0	1	0
kungens	king	0	0	1	0
kungens	the king's	0	0	1	0
svart	black	0	0	1	1
nyligen	recently	0	0	1	1
data	data	0	0	1	1
epost	e-mail	0	0	1	0
epost	email	0	0	1	0
portugisiska	portuguese	0	0	1	1
portugisiska	portugese	0	0	1	0
stress	stress	0	0	1	1
natural	natural	0	0	1	0
bergarter	rock types	0	0	1	0
bergarter	minerals	0	0	1	0
bergarter	rocks	0	0	1	0
undervisning	teaching	0	0	1	1
undervisning	undervising	0	0	1	0
undervisning	education	0	0	1	1
ss	ss	0	0	1	0
sr	sr	0	0	1	0
årlig	yearly	0	0	1	1
sv	sw	0	0	1	0
sv	south west	0	0	1	0
vikt	weight	0	0	1	1
st	saint	0	0	1	0
sk	so called	0	0	1	0
sk	known	0	0	1	0
so	so	0	0	1	0
sm	s-m	0	0	1	0
sm	swedish championship	0	0	1	0
sa	said	0	0	1	0
vika	fold	0	0	1	1
se	see	0	0	1	1
resulterar	resulting	0	0	1	0
resulterar	result	0	0	1	0
resulterar	results	0	0	1	0
allvarliga	serious	0	0	1	0
allvarliga	severe	0	0	1	0
resulterat	resulted	0	0	1	0
resulterat	resulted in	0	0	1	0
professorn	professor	0	0	1	0
professorn	the professor	0	0	1	0
kong	(hong) kong	0	0	1	0
kong	kong	0	0	1	0
antingen	presumably	0	0	1	0
antingen	either	0	0	1	1
förslaget	proposition	0	0	1	0
förslaget	the suggestion	0	0	1	0
förslaget	research team	0	0	1	0
upprätthåller	maintains	0	0	1	0
upprätthåller	maintaining	0	0	1	0
allvarligt	serious	0	0	1	0
allvarligt	severe	0	0	1	0
clinton	clinton	0	0	1	0
ingår	is	0	0	1	0
ingår	penetrations	0	0	1	0
torg	square	0	0	1	1
ingvar	ingvar	0	0	1	0
dialekter	dialects	0	0	1	0
människa	human being	0	0	1	0
människa	human	0	0	1	0
människa	man	0	0	1	1
torn	tower	0	0	1	1
tilldelats	assigned	0	0	1	0
tilldelats	awarded	0	0	1	0
turnera	tour	0	0	1	1
museu	museum	0	0	1	0
faderns	his father	0	0	1	0
faderns	the father's	0	0	1	0
monopol	monopoly	0	0	1	1
personlig	personal	0	0	1	1
svärd	sword	0	0	1	1
britter	britons	0	0	1	0
fastställa	determine	0	0	1	1
fastställa	confirm	0	0	1	0
konstnären	artist	0	0	1	0
konstnären	the artist	0	0	1	0
konstnären	artists	0	0	1	0
musiken	the music	0	0	1	0
musiken	music	0	0	1	0
matcher	matches	0	0	1	0
matcher	games	0	0	1	0
datorspel	video game	0	0	1	0
datorspel	computer game	0	0	1	0
nation	nation	0	0	1	1
records	records	0	0	1	0
förmågor	abilites	0	0	1	0
förmågor	capacities	0	0	1	0
förmågor	abilities	0	0	1	0
matchen	the game	0	0	1	0
matchen	match	0	0	1	0
kantoner	cantons	0	0	1	0
konstnärer	artists	0	0	1	0
musiker	musicians	0	0	1	0
musiker	musicants	0	0	1	0
lockar	attracts	0	0	1	0
lockar	curls	0	0	1	0
långbåge	longbow	1	1	0	0
långbåge	long arc	1	0	1	0
långbåge	many	1	0	1	0
långbåge	long bow	1	1	0	0
långbåge	ships	1	0	1	0
långbåge	angbage	1	0	1	0
långbåge	but spelt incorrectly below.	1	0	1	0
långbåge	i think it is language	1	0	1	0
långbåge	langbage	1	1	0	0
hjärtat	heart	0	0	1	0
hjärtat	the heart	0	0	1	0
sidor	pages	0	0	1	0
sidor	sides	0	0	1	0
sättas	turn	0	0	1	0
sättas	added	0	0	1	0
sättas	atta	0	0	1	0
dominerar	dominate	0	0	1	0
dominerar	dominates	0	0	1	0
domineras	dominated	0	0	1	0
runstenar	runestones	0	0	1	0
runstenar	rune stones	0	0	1	0
dominerat	docminaret	0	0	1	0
dominerat	dominated	0	0	1	0
föreställa	imagine	0	0	1	0
föreställa	pretend; imagine	0	0	1	0
prisma	prism	0	0	1	1
prisma	prisma	0	0	1	0
dynamiska	dynamic	0	0	1	0
greker	greek	0	0	1	0
greker	greeks	0	0	1	0
café	cafe	0	0	1	0
café	coffeehouse	0	0	1	0
café	café	0	0	1	0
delstaterna	states	0	0	1	0
jämna	even	0	0	1	0
hinduer	hindu	0	0	1	0
hinduer	hindus	0	0	1	0
krav	requirement	0	0	1	1
krav	conditions	0	0	1	0
krav	demands	0	0	1	0
riktigt	real	0	0	1	1
riktigt	right	0	0	1	0
ockupationen	the occupation	0	0	1	0
ockupationen	occupation	0	0	1	0
befolkningstillväxt	population growth	0	0	1	1
befolkningstillväxt	befolkningstillvaxt	0	0	1	0
måleri	painting	0	0	1	1
sjuka	disease	0	0	1	0
sjuka	sick	0	0	1	0
densitet	density	0	0	1	1
äga	be	0	0	1	0
äga	own	0	0	1	1
äga	aga	0	0	1	0
riktiga	real	0	0	1	0
internet	internet	0	0	1	0
roterar	rotates	0	0	1	0
bla	blah	0	0	1	0
bla	among others	0	0	1	0
arterna	the species	0	0	1	0
arterna	species	0	0	1	0
garantera	ensure	0	0	1	1
garantera	guarantee	0	0	1	1
singlar	singles	0	0	1	0
bytt	changed	0	0	1	0
bytt	traded	0	0	1	0
bytt	switched	0	0	1	0
byts	changed	0	0	1	0
byts	replaced	0	0	1	0
pilatus	pilatus	0	0	1	0
pilatus	pilate	0	0	1	1
osäker	insecure	0	0	1	1
osäker	unsure	0	0	1	1
byte	change of	0	0	1	0
byte	bytes	0	0	1	0
byta	switch	0	0	1	0
byta	change	0	0	1	1
byta	trade	0	0	1	1
sedd	seen	0	0	1	0
pund	pound	0	0	1	1
artister	artists	0	0	1	0
artister	performers	0	0	1	0
punk	punk rock	0	0	1	0
punk	punk	0	0	1	0
punk	para	0	0	1	0
flandern	flanders	0	0	1	1
dömande	sentencing	0	0	1	0
dömande	judging	0	0	1	0
massiva	solid	0	0	1	0
massiva	massive	0	0	1	0
artisten	the artist	0	0	1	0
artisten	artist	0	0	1	0
gordon	gordon	0	0	1	0
givits	given	0	0	1	0
följt	followed	0	0	1	0
förutom	apart from	0	0	1	0
förutom	besides; in addition to; aside from	0	0	1	0
förutom	except	0	0	1	0
väpnad	armed	0	0	1	1
potter	potter	0	0	1	0
potter	pots	0	0	1	0
one	one	0	0	1	0
tsunamier	tsunamis	0	0	1	0
bekräftades	confirmed	0	0	1	0
bekräftades	was confirmed	0	0	1	0
open	open	0	0	1	1
ont	bad	0	0	1	0
urin	urine	0	0	1	1
city	city	0	0	1	0
tekniska	technical	0	0	1	0
uppnådde	met	0	0	1	0
uppnådde	achieved	0	0	1	0
flytande	floating	0	0	1	1
flytande	liquid	0	0	1	1
teologi	teology	0	0	1	0
teologi	theology	0	0	1	1
gasen	gas	0	0	1	0
intill	beside	0	0	1	0
intill	adjacent to	0	0	1	0
intill	adjacent	0	0	1	1
williams	williams	0	0	1	0
animerade	animated	0	0	1	1
vilka	who; which; that	0	0	1	0
vilka	who	0	0	1	1
vilka	which	0	0	1	1
£m	million pounds	0	0	1	0
löfte	promise	0	0	1	1
bär	carryng	0	0	1	0
bär	here	0	0	1	0
bär	berries	0	0	1	0
irakiska	iraqi	0	0	1	0
irakiska	irakish	0	0	1	0
svenskarna	the swedes	0	0	1	0
svenskarna	swedes	0	0	1	0
synsättet	approach	0	0	1	0
synsättet	view	0	0	1	0
yttersta	furthest	0	0	1	0
yttersta	supreme	0	0	1	0
yttersta	highly	0	0	1	0
provins	province	0	0	1	1
dygn	day	0	0	1	1
fiskar	fishes	0	0	1	0
fiskar	fish	0	0	1	0
uppenbarelser	revelations	0	0	1	0
berlinmuren	berlin wall	0	0	1	0
berlinmuren	the berlin wall	0	0	1	0
föreslagit	suggested	0	0	1	0
föreslagit	proposed	0	0	1	0
uppfördes	was constructed	0	0	1	0
uppfördes	built	0	0	1	0
uppfördes	constructed	0	0	1	0
kamprad	kamprad	0	0	1	0
tankar	tank	0	0	1	0
tankar	thoughts	0	0	1	0
sak	thing	0	0	1	1
sak	matter; case	0	0	1	0
sak	substance	0	0	1	0
san	san	0	0	1	0
sam	co	0	0	1	0
generation	generation	0	0	1	0
konsekvenser	consequences	0	0	1	0
argument	argument	0	0	1	1
argument	arguments	0	0	1	0
överhuvudtaget	in general	0	0	1	0
överhuvudtaget	generally	0	0	1	0
överhuvudtaget	on the whole	0	0	1	1
burundi	burundi	0	0	1	0
allen	allen	0	0	1	0
turner	tournament	0	0	1	0
staden	city	0	0	1	0
staden	the city	0	0	1	0
priserna	prices	0	0	1	0
priserna	the prices	0	0	1	0
indelad	divided	0	0	1	0
skickades	was sent	0	0	1	0
skickades	sent	0	0	1	0
takt	rate	0	0	1	1
zon	zone	0	0	1	1
zoo	zoo	0	0	1	1
jefferson	jefferson	0	0	1	0
massa	mass	0	0	1	1
begreppen	the concepts	0	0	1	0
begreppen	the terms	0	0	1	0
begreppen	terms	0	0	1	0
muslimer	mulismer	0	0	1	0
muslimer	muslims	0	0	1	0
plattform	lost	1	0	1	0
plattform	stage; platform	1	0	1	0
plattform	platform; stand	1	0	1	0
plattform	platform	1	1	1	1
plattform	pad	1	1	1	0
plattform	stand	1	0	1	0
plattform	the plates	1	0	1	0
plattform	rig	1	1	0	0
plattform	old plate	1	0	1	0
plattform	plattform	1	0	1	0
finlands	finland's	0	0	1	0
finlands	finlands	0	0	1	0
sekreterare	secretary	0	0	1	1
därpå	then	0	0	1	1
därpå	thereon	0	0	1	1
därpå	darpa	0	0	1	0
mynt	coins	0	0	1	0
mynt	coin	0	0	1	1
religionen	religion	0	0	1	0
religionen	the religion	0	0	1	0
pastor	pastor	0	0	1	1
religioner	religions	0	0	1	0
forskningen	the science	0	0	1	0
forskningen	research	0	0	1	0
översikt	overview	0	0	1	1
översikt	over term	0	0	1	0
beväpnade	armed	0	0	1	0
kontroversiell	controversial herring	0	0	1	0
kontroversiell	controversial	0	0	1	1
höjd	height; above	0	0	1	0
höjd	height	0	0	1	1
höja	increase	0	0	1	0
höja	hoja	0	0	1	0
höja	raise	0	0	1	1
driva	operate	0	0	1	1
driva	run	0	0	1	0
phil	phil	0	0	1	0
inledningen	introduction	0	0	1	0
inledningen	the beginning	0	0	1	0
inledningen	the introduction	0	0	1	0
ursprung	origin	0	0	1	1
ursprung	root	0	0	1	1
fredspriset	nobel peace prize	0	0	1	0
fredspriset	peace price	0	0	1	0
fredspriset	peace prize	0	0	1	0
rykte	reputation	0	0	1	1
sades	said	0	0	1	0
sades	was said	0	0	1	0
katekes	catechism	0	0	1	1
engagemang	commitment	0	0	1	1
olagligt	illegal	0	0	1	0
axl	axl	0	0	1	0
beckham	beckham	0	0	1	0
dimensioner	dimensions	0	0	1	0
klimatologi	use	1	0	1	0
klimatologi	klimatology	1	0	1	0
klimatologi	klimatologia	1	1	0	0
klimatologi	climateology	1	0	1	0
klimatologi	have	1	0	1	0
klimatologi	climatology	1	1	0	0
börja	start	0	0	1	1
börje	borje	0	0	1	0
börje	börje	0	0	1	0
antalet	number	0	0	1	0
antalet	the number	0	0	1	0
föreningen	the association	0	0	1	0
föreningen	association	0	0	1	0
föreningen	compound	0	0	1	0
slog	hit	0	0	1	0
hockey	ice hockey	0	0	1	1
hockey	hockey	0	0	1	1
caroline	caroline	0	0	1	0
carolina	carolina	0	0	1	0
beatles	beatles	0	0	1	0
kategorimusik	category music	0	0	1	0
fader	father	0	0	1	1
populär	popular	0	0	1	1
berör	affecting	0	0	1	0
berör	affect	0	0	1	0
berör	concerns	0	0	1	0
avrättningar	execution	0	0	1	0
avrättningar	executions	0	0	1	0
härrör	derived	0	0	1	0
platta	flat	0	0	1	1
spetshundar	sets dogs	0	0	1	0
spetshundar	tip of dogs	0	0	1	0
artist	artist	0	0	1	1
roger	roger	0	0	1	0
ljudet	the sound	0	0	1	0
ljudet	noise	0	0	1	0
varna	varna	0	0	1	0
varna	alerting	0	0	1	0
monark	monarch	0	0	1	1
vision	vision	0	0	1	1
spetsen	edge; top	0	0	1	0
spetsen	tip	0	0	1	0
snabbare	rapid	0	0	1	0
snabbare	faster	0	0	1	0
uppnått	met	0	0	1	0
uppnått	achieved	0	0	1	0
behovet	need	0	0	1	0
behovet	the need	0	0	1	0
up	i[	0	0	1	0
up	up	0	0	1	0
värre	worse	0	0	1	1
talman	spokesperson	0	0	1	0
talman	president	0	0	1	0
talman	speaker	0	0	1	1
enhetlig	single	0	0	1	0
enhetlig	unitary	0	0	1	1
enhetlig	uniform	0	0	1	1
kritiserade	critisized	0	0	1	0
kritiserade	criticized	0	0	1	0
kritiserade	criticised	0	0	1	0
upplever	experiencing	0	0	1	0
upplever	experience	0	0	1	0
kontrakt	agreement	0	0	1	1
kontrakt	contract	0	0	1	1
kilometer	kilometer	0	0	1	1
kilometer	kilometers	0	0	1	0
färgerna	colors	0	0	1	0
amerikanskt	american	0	0	1	0
utföras	be	0	0	1	0
utföras	performed	0	0	1	0
anledningarna	reasons	0	0	1	0
anledningarna	the reasons	0	0	1	0
screen	screen	0	0	1	0
fynd	finding; finds	0	0	1	0
fynd	findings	0	0	1	0
upphovsrätt	rise knob	0	0	1	0
upphovsrätt	copyright	0	0	1	1
pågick	manufacture was	0	0	1	0
pågick	lasted	0	0	1	0
amerikanske	american	0	0	1	0
amerikanske	the american	0	0	1	0
awards	awards	0	0	1	0
jobb	job	0	0	1	1
jobb	work	0	0	1	1
amerikanska	u.s.	0	0	1	0
amerikanska	american	0	0	1	0
mariette	mariette	0	0	1	0
basisten	basist	0	0	1	0
basisten	bassist	0	0	1	0
basisten	the basist	0	0	1	0
skär	will	0	0	1	0
skär	cut	0	0	1	0
skär	skerry	0	0	1	1
mans	man's	0	0	1	0
föras	be	0	0	1	0
föras	be brought	0	0	1	0
föras	taken to	0	0	1	0
rädsla	fear	0	0	1	1
s	s	0	0	1	0
hälsa	health	0	0	1	1
hälsa	tell (him i said hi)	0	0	1	0
hälsa	neck	0	0	1	0
mani	mani	0	0	1	0
mani	mania	0	0	1	1
skäl	reasons	0	0	1	0
skäl	reason	0	0	1	1
härstamma	originate	0	0	1	1
härstamma	stem	0	0	1	0
upproret	the upprising	0	0	1	0
upproret	revolt	0	0	1	0
upproret	rebellion	0	0	1	0
klimat	climate	0	0	1	1
hamnade	landed	0	0	1	0
hamnade	ended up	0	0	1	0
anta	assume	0	0	1	0
anta	adopting	0	0	1	0
anta	assume; adopt	0	0	1	0
samtal	call	0	0	1	1
samtal	conersation	0	0	1	0
drogs	was pulled	0	0	1	0
drogs	was	0	0	1	0
främre	forward	0	0	1	1
främre	front	0	0	1	1
främre	anterior	0	0	1	1
teddy	teddy	0	0	1	0
farfar	paternal grandfather	0	0	1	0
farfar	grandfather	0	0	1	1
west	west	0	0	1	0
airlines	airlines	0	0	1	0
bolag	company	0	0	1	1
luft	air	0	0	1	1
cupen	the cup	0	0	1	0
cupen	cup	0	0	1	0
lidit	sustained	0	0	1	0
lidit	suffered	0	0	1	0
vänner	friendas	0	0	1	0
vänner	friends	0	0	1	0
formen	the form	0	0	1	0
formen	form	0	0	1	0
formel	formula	0	0	1	1
arabiska	arabic	0	0	1	1
arabiska	arabian	0	0	1	0
diktaturen	dictatorship	0	0	1	0
warhol	warhol	0	0	1	0
former	forms	0	0	1	0
landskapen	the landscapes	0	0	1	0
landskapen	landscapes	0	0	1	0
landskapen	landscape	0	0	1	0
samling	concentration	0	0	1	0
samling	collection	0	0	1	1
mona	mona	0	0	1	0
landskapet	landscape	0	0	1	0
norrköpings	norrköpings	0	0	1	0
situation	situation	0	0	1	1
situation	position	0	0	1	0
återfanns	was rediscovered	0	0	1	0
återfanns	found	0	0	1	0
återfanns	can be found	0	0	1	0
peruanska	peruvian	0	0	1	0
peruanska	peruan	0	0	1	0
förlorar	loss	0	0	1	0
förlorar	loses	0	0	1	0
ive	i've	0	0	1	0
aluminium	aluminum	0	0	1	1
förlorat	lost	0	0	1	0
startar	begins	0	0	1	0
startar	start	0	0	1	0
startar	starts	0	0	1	0
bror	brother	0	0	1	1
bron	bridge	0	0	1	0
bron	the bridge	0	0	1	0
jenny	jenny	0	0	1	0
bestämmelser	regulations	0	0	1	0
bestämmelser	measures	0	0	1	0
bestämmelser	conditions	0	0	1	0
sammanfaller	coinciding	0	0	1	0
sammanfaller	coincides	0	0	1	0
omnämns	mentioned	0	0	1	0
omnämns	is mentioned	0	0	1	0
hästens	horses	0	0	1	0
hästens	horse's	0	0	1	0
hästens	horse	0	0	1	0
linje	line	0	0	1	1
wilhelm	wilhelm	0	0	1	0
otto	otto	0	0	1	0
oceanen	the ocean	0	0	1	0
oceanen	ocean	0	0	1	0
hämta	retrieve	0	0	1	0
hämta	fetch	0	0	1	1
ekologi	ecology	0	0	1	1
ludwig	lugwig	0	0	1	0
ludwig	ludwig	0	0	1	0
nationalparker	national parks	0	0	1	0
värmestrålningen	heat radiation	0	0	1	0
singapore	singapore	0	0	1	0
fåglar	birds	0	0	1	0
lindgrens	lindgren's	0	0	1	0
lindgrens	lindgrens	0	0	1	0
lindgrens	lindgren	0	0	1	0
cullen	cullen	0	0	1	0
senator	senator	0	0	1	1
dsmiv	dsm-iv	0	0	1	0
försvarare	defenders	0	0	1	0
försvarare	defender	0	0	1	1
costa	costa	0	0	1	0
rorsman	rosman	1	0	1	0
rorsman	steersman	1	1	0	1
rorsman	helms man	1	0	1	0
rorsman	usage	1	0	1	0
rorsman	using	1	0	1	0
rorsman	helmsman	1	1	0	1
avser	regard	0	0	1	0
avser	regards	0	0	1	0
avser	refers to	0	0	1	0
avses	refered	0	0	1	0
avses	regard	0	0	1	0
avses	referred	0	0	1	0
iraks	iraq	0	0	1	0
gudomliga	gudombliga	0	0	1	0
gudomliga	divine	0	0	1	0
summer	sommar	0	0	1	0
edwards	edwards	0	0	1	0
edwards	edward's	0	0	1	0
uppmärksammade	observed	0	0	1	0
uppmärksammade	noted	0	0	1	0
uppmärksammade	noticed	0	0	1	0
igelkottar	hedgehogs	0	0	1	0
tätorter	urban	0	0	1	0
tätorter	conurbation	0	0	1	0
tätorter	cities	0	0	1	0
rest	remain	0	0	1	0
rest	residual	0	0	1	1
rest	rest	0	0	1	1
tätorten	conurbation	0	0	1	0
tätorten	agglomeration	0	0	1	0
bergman	bergman	0	0	1	0
koncentration	concentration	0	0	1	1
utnyttja	use	0	0	1	1
psykologisk	psychological	0	0	1	1
likheter	similarities	0	0	1	0
likheter	similarity	0	0	1	0
resa	travel	0	0	1	1
libyen	libya	0	0	1	1
judarnas	jews	0	0	1	0
kastar	castes	0	0	1	0
kastar	throws	0	0	1	0
kastar	to throw	0	0	1	0
avgå	resign	0	0	1	1
heliga	saints	0	0	1	0
heliga	holy	0	0	1	0
heliga	holy; holy	0	0	1	0
unika	unique	0	0	1	0
sprider	spread	0	0	1	0
sprider	spreads out	0	0	1	0
sprider	spreads	0	0	1	0
armén	the army	0	0	1	0
helige	holy	0	0	1	0
låtskrivare	songwriter	0	0	1	0
låtskrivare	song writers	0	0	1	0
instrument	intrument	0	0	1	0
får	may be	0	0	1	0
får	can	0	0	1	0
får	allow	0	0	1	0
växte	grew	0	0	1	0
växte	grow	0	0	1	0
unikt	unique	0	0	1	0
heligt	holy	0	0	1	0
heligt	heligit	0	0	1	0
riksväg	national highway	0	0	1	0
riksväg	highway	0	0	1	0
tjänare	servant	0	0	1	1
motorvägar	highways	0	0	1	0
motorvägar	motor	0	0	1	0
snart	soon	0	0	1	1
snart	once	0	0	1	0
huvudvärk	headache	0	0	1	1
återkom	return	0	0	1	0
återkom	returned	0	0	1	0
återkom	feedback	0	0	1	0
vinkel	angle	0	0	1	1
dark	dark	0	0	1	0
regim	regimen	0	0	1	1
regim	regime	0	0	1	1
unesco	unesco	0	0	1	0
skadade	wounded	0	0	1	0
skadade	damaged	0	0	1	0
stammar	strains	0	0	1	0
stammar	stutters	0	0	1	0
stammar	tribes	0	0	1	0
statsreligion	state religion	0	0	1	0
bekräftar	confirmed	0	0	1	0
bekräftar	confirms	0	0	1	0
bekräftar	confirming	0	0	1	0
framsteg	progress	0	0	1	1
bekräftat	confirmed	0	0	1	0
träda	esterified	0	0	1	0
träda	emerge	0	0	1	0
träda	fallow	0	0	1	1
tvserie	tv serial	0	0	1	0
tsunami	tsunami	0	0	1	0
ekonomier	economies	0	0	1	0
stupade	fallen	0	0	1	0
stupade	killed	0	0	1	0
fossila	fossilized	0	0	1	0
fossila	fossil	0	0	1	0
inter	inter	0	0	1	0
intet	nothing	0	0	1	1
intet	no	0	0	1	0
magnetfält	magnetic	0	0	1	0
magnetfält	magnetic field	0	0	1	1
brita	brita	0	0	1	0
domkyrkan	cathedral	0	0	1	0
domkyrkan	the cathedral	0	0	1	0
älgar	moose	0	0	1	0
ursprungsbefolkning	native population	0	0	1	0
ursprungsbefolkning	indigenous	0	0	1	0
märke	badge	0	0	1	0
märke	label	0	0	1	1
ekman	ekman	0	0	1	0
försvinner	disappears	0	0	1	0
försvinner	disappearing	0	0	1	0
försvinner	disappear	0	0	1	0
märks	notice	0	0	1	0
märks	labeled	0	0	1	0
märks	noted	0	0	1	0
strindberg	strindberg	0	0	1	0
institutionerna	institutions	0	0	1	0
företaget	the company	0	0	1	0
ddr	ddr	0	0	1	0
exil	exile	0	0	1	1
cannabis	cannabis	0	0	1	1
miljö	environment	0	0	1	1
företagen	the companies	0	0	1	0
företagen	taken present	0	0	1	0
katolsk	catholic	0	0	1	1
stränder	beaches	0	0	1	0
jacksons	jackson's	0	0	1	0
jacksons	jacksons	0	0	1	0
jacksons	jackson	0	0	1	0
medlemsstater	member	0	0	1	0
medlemsstater	member states	0	0	1	0
medlemsstater	member-state	0	0	1	0
påverka	impact	0	0	1	0
påverka	influence	0	0	1	1
stone	least	0	0	1	0
organisationen	organization	0	0	1	0
organisationen	the organization	0	0	1	0
ace	ace	0	0	1	0
herrlandslag	men's national team	0	0	1	0
herrlandslag	women's national teams	0	0	1	0
andreas	andreas	0	0	1	0
vissa	some	0	0	1	0
populationen	the population	0	0	1	0
populationen	population	0	0	1	0
befinner	is	0	0	1	0
befinner	placed; situated; positioned; are	0	0	1	0
populationer	populations	0	0	1	0
wien	vienna	0	0	1	1
organisationer	organizations	0	0	1	0
organisationer	organisations	0	0	1	0
industri	industry	0	0	1	1
industri	industrial	0	0	1	0
bond	bond	0	0	1	0
visst	specific	0	0	1	0
visst	certain	0	0	1	0
billboardlistan	billboard list	0	0	1	0
billboardlistan	bilboardlist	0	0	1	0
berger	berger	0	0	1	0
upplevelser	experiences	0	0	1	0
ronden	round	0	0	1	0
bryts	breaks	0	0	1	0
nationalencyklopedin	national encyclopedia	0	0	1	0
nationalencyklopedin	the national encyclopedia	0	0	1	0
image	image	0	0	1	1
partiet	the party	0	0	1	0
partiet	portion	0	0	1	0
bryta	break	0	0	1	1
partier	portions	0	0	1	0
partier	parties	0	0	1	0
bergen	the mountains	0	0	1	0
bergen	mountain	0	0	1	0
bergen	mountains	0	0	1	0
het	hot	0	0	1	1
het	up to date	0	0	1	0
utövade	exerted	0	0	1	0
utövade	exercised	0	0	1	0
kategorifödda	category born	0	0	1	0
kategorifödda	category: born	0	0	1	0
kallats	was called	0	0	1	0
kallats	called	0	0	1	0
philadelphia	philadelphia	0	0	1	0
evangeliska	evangelical	0	0	1	0
legitimitet	legitimacy	0	0	1	1
förmåga	abilities	0	0	1	0
förmåga	ability	0	0	1	1
hel	full	0	0	1	1
hel	(whole) lot (of)	0	0	1	0
hem	home	0	0	1	1
hem	dobladillo	0	0	1	0
hem	back	0	0	1	0
hamnen	harbour	0	0	1	0
hamnen	the harbour	0	0	1	0
sover	sleep	0	0	1	0
enorm	huge	0	0	1	1
enorm	enormous	0	0	1	1
dagen	day	0	0	1	0
complete	complete	0	0	1	0
norrköping	norrköping	0	0	1	0
bevarat	preserve	0	0	1	0
bevarat	preserved	0	0	1	0
bevaras	are protected	0	0	1	0
bevaras	preserved	0	0	1	0
mick	microphone	0	0	1	0
mick	mick	0	0	1	0
mick	mike (microphone)	0	0	1	0
kontroverser	controversies	0	0	1	0
kontroverser	contraversies	0	0	1	0
existerande	current	0	0	1	0
existerande	existing	0	0	1	1
bevarad	kept	0	0	1	0
bevarad	preserved	0	0	1	1
störta	rush	0	0	1	0
störta	crash	0	0	1	0
störta	interfere	0	0	1	0
jamaicas	jamaicas	0	0	1	0
jamaicas	jamaica's	0	0	1	0
hexadecimalt	hexa-decimal	0	0	1	0
hexadecimalt	hex	0	0	1	0
kvartsfinalen	quarter finals	0	0	1	0
kvartsfinalen	quarterfinals	0	0	1	0
vinkeln	angle	0	0	1	0
vinkeln	the angle	0	0	1	0
afrodite	aphrodite	0	0	1	0
afrodite	afrodite	0	0	1	0
karriär	career	0	0	1	1
age	do	0	0	1	0
age	age	0	0	1	0
puls	pulse	0	0	1	1
ac	ac	0	0	1	0
ab	ab	0	0	1	0
brodern	the brother	0	0	1	0
brodern	brother	0	0	1	0
johnny	johny	0	0	1	0
johnny	johnny	0	0	1	0
redovisas	reported	0	0	1	0
redovisas	shown	0	0	1	0
redovisas	accounted for	0	0	1	0
gustafs	gustafs	0	0	1	0
gustafs	gustaf's	0	0	1	0
am	am	0	0	1	0
al	alder	0	0	1	1
an	an	0	0	1	0
as	as	0	0	1	1
beordrade	commanded	0	0	1	0
beordrade	ordered	0	0	1	0
au	au	0	0	1	0
at	at	0	0	1	0
av	of	0	0	1	1
testamentet	testament	0	0	1	0
vore	would	0	0	1	0
vore	were	0	0	1	0
federala	federal	0	0	1	0
axelmakterna	the axis	0	0	1	0
axelmakterna	axis	0	0	1	0
premiär	prime	0	0	1	0
premiär	premiere	0	0	1	1
sköter	handles	0	0	1	0
sköter	handle	0	0	1	0
gifta	marry	0	0	1	0
gifta	married	0	0	1	0
koppar	copper	0	0	1	1
gifte	married	0	0	1	0
medverkan	the contribution	0	0	1	0
medverkan	participation	0	0	1	1
kvarstod	remained	0	0	1	0
öland	oland	0	0	1	0
öland	öland	0	0	1	0
terra	terra	0	0	1	1
medverkat	participated	0	0	1	0
medverkar	contribute	0	0	1	0
medverkar	contributes	0	0	1	0
förälskad	in love	0	0	1	1
terry	terry	0	0	1	0
ekonomi	economic	0	0	1	0
ekonomi	economy	0	0	1	1
dokumentär	documentary	0	0	1	1
forntida	pristine	0	0	1	1
forntida	ancient	0	0	1	1
forntida	prehistoric	0	0	1	0
kommunen	municipality	0	0	1	0
kommuner	municipalities	0	0	1	0
kommuner	local	0	0	1	0
kommuner	counties	0	0	1	0
beteckning	indication	0	0	1	1
beteckning	label	0	0	1	0
adam	adam	0	0	1	0
omgivningen	surroundings	0	0	1	0
omgivningen	the surrounding	0	0	1	0
omgivningen	ambient	0	0	1	0
hjälp	using	0	0	1	0
hjälp	help	0	0	1	1
original	original	0	0	1	1
original	orignal	0	0	1	0
islamiska	islamic	0	0	1	0
resor	travels	0	0	1	0
resor	travel	0	0	1	0
elektron	electron	0	0	1	1
halsen	throat	0	0	1	0
halsen	the neck	0	0	1	0
halsen	the throat	0	0	1	0
anpassning	adaption	0	0	1	0
anpassning	adjustment	0	0	1	1
kammare	chamber	0	0	1	1
likartade	similiar	0	0	1	0
likartade	similar	0	0	1	0
avslöjade	revealed	0	0	1	0
reduktion	reduction	1	1	0	0
reduktion	processes	1	0	1	0
norr	north	0	0	1	1
skogarna	the forests	0	0	1	0
skogarna	forests	0	0	1	0
störning	noise	0	0	1	0
störning	high accession	0	0	1	0
ullevi	ullevi	0	0	1	0
tv	tv	0	0	1	1
romanen	novel	0	0	1	0
to	to	0	0	1	0
mildare	cooler	0	0	1	0
mildare	milder	0	0	1	0
mildare	mild	0	0	1	0
romaner	novels	0	0	1	0
th	th	0	0	1	0
nord	north	0	0	1	1
gör	does	0	0	1	0
gör	makes	0	0	1	0
te	tea	0	0	1	1
östafrika	east africa	0	0	1	0
ta	to	0	0	1	0
ta	take	0	0	1	1
ghana	ghana	0	0	1	1
hämtat	collected	0	0	1	0
hämtat	downloaded	0	0	1	0
hämtat	taken	0	0	1	0
händelserna	the events	0	0	1	0
händelserna	events	0	0	1	0
händelserna	the happenings	0	0	1	0
arvet	the inheritance	0	0	1	0
arvet	heritage	0	0	1	0
telefonen	phone	0	0	1	0
telefonen	the telephone	0	0	1	0
strand	beach	0	0	1	1
sant	true	0	0	1	0
ensamma	alone	0	0	1	0
djurarter	species of animals	0	0	1	0
djurarter	animal species	0	0	1	0
djurarter	species	0	0	1	0
borrelia	borrelia	0	0	1	0
borrelia	borreliosis	0	0	1	0
venezuela	venezuela	0	0	1	0
utvisning	penalty	0	0	1	0
utvisning	expulsion	0	0	1	0
muslimska	muslim	0	0	1	0
sand	sand	0	0	1	1
sand	sandy	0	0	1	0
siffrorna	the numbers	0	0	1	0
siffrorna	figures	0	0	1	0
siffrorna	numbers	0	0	1	0
smala	narrow	0	0	1	0
harry	harry	0	0	1	0
sann	true	0	0	1	1
samoa	samoa	0	0	1	0
rapporter	reports	0	0	1	0
synd	sin	0	0	1	1
rörde	had something to do with	0	0	1	0
rörde	touched	0	0	1	0
rörde	was about	0	0	1	0
skede	period	0	0	1	1
skede	analysis	0	0	1	0
skede	stage	0	0	1	0
påbörjades	commenced; begun	0	0	1	0
påbörjades	initiated	0	0	1	0
påbörjades	was started	0	0	1	0
givaren	donor	0	0	1	0
givaren	the giver	0	0	1	0
givaren	dealer	0	0	1	0
brottet	offense	0	0	1	0
brottet	the crime	0	0	1	0
brottet	the crime; offense; infraction; transgression	0	0	1	0
syns	seen	0	0	1	0
syns	visible	0	0	1	0
richard	richard	0	0	1	0
stjäla	steal	0	0	1	1
stjäla	stealing	0	0	1	0
övrig	other	0	0	1	1
soldater	soldiers	0	0	1	0
islams	islams	0	0	1	0
islams	islam's	0	0	1	0
leif	leif	0	0	1	0
gjorts	made	0	0	1	0
gjorts	done	0	0	1	0
full	full	0	0	1	1
gruppen	the group	0	0	1	0
gruppen	group	0	0	1	0
människors	humans	0	0	1	0
människors	human	0	0	1	0
människors	people's	0	0	1	1
arkeologiska	archaeological	0	0	1	0
november	november	0	0	1	1
legend	legend	0	0	1	1
sålda	sold	0	0	1	0
sålda	salda	0	0	1	0
sålde	sold	0	0	1	0
sålde	sells drinks	0	0	1	0
kräva	require	0	0	1	0
kräva	demand	0	0	1	1
inverkan	impact	0	0	1	1
inverkan	influence	0	0	1	1
inverkan	effect	0	0	1	0
exklusiv	exclusive	0	0	1	1
krävt	taken	0	0	1	0
krävt	required	0	0	1	0
krävs	needs	0	0	1	0
krävs	required	0	0	1	0
krävs	requires	0	0	1	0
social	social	0	0	1	1
action	action	0	0	1	0
oftare	more	0	0	1	0
oftare	more often	0	0	1	0
oftare	more frequently	0	0	1	0
varelser	creatures	0	0	1	0
hamnar	lands	0	0	1	0
hamnar	ports	0	0	1	0
kommunistpartiet	communist party	0	0	1	0
kommunistpartiet	the communist party	0	0	1	0
vid	by	0	0	1	1
vid	at	0	0	1	1
vid	in	0	0	1	0
ordinarie	ordinary	0	0	1	1
ordinarie	permanent	0	0	1	1
ordinarie	regular	0	0	1	0
vii	vii	0	0	1	0
vin	whine	0	0	1	0
vin	wine	0	0	1	1
hamnat	got	0	0	1	0
hamnat	ended up	0	0	1	0
hamnat	got in to	0	0	1	0
juridiskt	legally	0	0	1	0
juridiskt	juridical	0	0	1	0
juridiskt	judicial	0	0	1	0
vis	vis	0	0	1	0
vis	wise	0	0	1	1
vis	way	0	0	1	1
vit	white	0	0	1	1
spelaren	the player	0	0	1	0
skapa	create	0	0	1	1
skapa	creating	0	0	1	0
skapa	bushel	0	0	1	0
biskopen	bishop	0	0	1	0
biskopen	the bishop	0	0	1	0
bränslen	fuel	0	0	1	0
bränslen	fuels	0	0	1	0
klädsel	cover	0	0	1	0
strömningar	tendencies	0	0	1	0
strömningar	sentiments	0	0	1	0
mors	mothers	0	0	1	0
mors	mother	0	0	1	0
petroleum	oil	0	0	1	0
petroleum	petroleum	0	0	1	1
underordnade	subordinate	0	0	1	0
underordnade	subordinates	0	0	1	0
pearl	pearl	0	0	1	0
sitter	is	0	0	1	0
sitter	serve	0	0	1	0
sitter	sit	0	0	1	0
presenterades	presented	0	0	1	0
rhen	the rhine	0	0	1	0
rhen	rhine	0	0	1	1
öka	oka	0	0	1	0
öka	increase	0	0	1	1
öka	increasing	0	0	1	0
mora	mora	0	0	1	0
bevis	certificate	0	0	1	1
bevis	evidence	0	0	1	1
mord	murder	0	0	1	1
ragnar	ragnar	0	0	1	0
uppskattad	estimated	0	0	1	0
uppskattad	appreciated	0	0	1	0
ögonen	eyes	0	0	1	0
ögonen	the eyes	0	0	1	0
uppskattas	is appreciated	0	0	1	0
uppskattas	estimated	0	0	1	0
uppskattas	appreciated	0	0	1	0
uppskattar	estimated	0	0	1	0
uppskattar	estimates	0	0	1	0
schweiz	switzerland	0	0	1	1
socialt	socially	0	0	1	0
socialt	social	0	0	1	0
medelklassen	middle class	0	0	1	0
science	science	0	0	1	0
försvarsmakt	armed forces	0	0	1	0
faser	phase	0	0	1	0
faser	phases	0	0	1	0
dancehall	dance hall	0	0	1	0
dancehall	dancehall	0	0	1	0
omständigheter	event	0	0	1	0
omständigheter	circumstances	0	0	1	1
klp	klp	0	0	1	0
cykel	bicycle	0	0	1	1
cykel	cycle	0	0	1	1
morgan	morgan	0	0	1	0
kapitalism	capitalism	0	0	1	1
studenter	students	0	0	1	0
jakob	jakob	0	0	1	0
skadliga	harmful	0	0	1	0
skadliga	deleterious	0	0	1	0
våglängder	wavelength	0	0	1	0
våglängder	wave lengths	0	0	1	0
våglängder	wavelengths	0	0	1	0
staten	state	0	0	1	0
mellersta	middle	0	0	1	1
mellersta	the middle	0	0	1	0
states	states	0	0	1	0
stater	states	0	0	1	0
spansk	spanish	0	0	1	1
återkomst	return	0	0	1	1
information	information	0	0	1	1
hugo	hugo	0	0	1	0
uppfattade	perceived	0	0	1	0
uppfattade	perceive	0	0	1	0
förhandlingar	negotiations	0	0	1	0
läran	teaching	0	0	1	0
läran	the teaching	0	0	1	0
läran	laran	0	0	1	0
ansetts	considered	0	0	1	0
ansetts	regarded	0	0	1	0
ansetts	regarded; viewed (as)	0	0	1	0
världshälsoorganisationen	world health organization	0	0	1	0
lejon	lion	0	0	1	1
bröllop	brollop	0	0	1	0
bröllop	wedding	0	0	1	1
behöva	need	0	0	1	1
riksdagens	the parliament's	0	0	1	0
riksdagens	the parliaments	0	0	1	0
retorik	rhetoric	0	0	1	1
variant	type	0	0	1	0
variant	variant	0	0	1	1
variant	variety	0	0	1	0
långsamma	slow	0	0	1	0
kedjan	chain	0	0	1	0
kedjan	the chain	0	0	1	0
produktionen	production	0	0	1	0
produktionen	the production	0	0	1	0
användas	used	0	0	1	0
referens	reference	0	0	1	1
lanka	lanka	0	0	1	0
lanka	(sri) lanka	0	0	1	0
står	standing	0	0	1	0
står	star	0	0	1	0
står	stand	0	0	1	0
barnens	children's	0	0	1	0
barnens	the child's	0	0	1	0
barnens	childrens	0	0	1	0
komplext	complex	0	0	1	0
anklagade	accused	0	0	1	0
pucken	the puck	0	0	1	0
sjön	sjon	0	0	1	0
sjön	lake	0	0	1	0
förändras	fora preferred	0	0	1	0
förändras	changes	0	0	1	0
komplexa	complex	0	0	1	0
utvidgning	enlargement; expansion	0	0	1	0
utvidgning	enlargement	0	0	1	1
tål	can take	0	0	1	0
tål	stand	0	0	1	0
tål	is resistant to	0	0	1	0
nationerna	the nations	0	0	1	0
nationerna	nations	0	0	1	0
blommor	flowers	0	0	1	0
resurs	resusrs	1	0	1	0
resurs	resurs	1	0	1	0
resurs	resource	1	1	0	1
resurs	factory	1	0	1	0
resurs	resources	1	0	1	0
trade	esterified	0	0	1	0
scott	scott	0	0	1	0
kvinnors	women	0	0	1	0
kvinnors	women's	0	0	1	0
aktiviteter	activities	0	0	1	0
aktiviteter	activity	0	0	1	0
årig	year old	0	0	1	0
årig	minor	0	0	1	0
radion	the radio	0	0	1	0
radion	radio	0	0	1	0
vietnamkriget	the vietnam war	0	0	1	0
vietnamkriget	vietnam war	0	0	1	0
läses	read	0	0	1	0
läses	is read	0	0	1	0
läser	read	0	0	1	0
läser	are reading	0	0	1	0
behålla	container	0	0	1	0
behålla	keep	0	0	1	1
alla	all	0	0	1	1
alla	everyone	0	0	1	1
protestanter	protestants	0	0	1	0
caesars	caesars	0	0	1	0
termen	the term	0	0	1	0
termen	term	0	0	1	0
hounds	hounds	0	0	1	0
termer	term	0	0	1	0
termer	terms	0	0	1	0
allt	all	0	0	1	1
alls	all	0	0	1	0
stadshus	town hall	0	0	1	1
stadshus	city hall; town hall	0	0	1	0
isaac	isaac	0	0	1	0
isaac	issac	0	0	1	0
strålning	radiation	0	0	1	1
ungefär	approx.; approximately	0	0	1	0
ungefär	about	0	0	1	1
ungefär	approximately	0	0	1	1
krävdes	were required	0	0	1	0
privilegier	privileges	0	0	1	0
förespråkade	advocate	0	0	1	0
förespråkade	advocated	0	0	1	0
inledande	initial	0	0	1	1
produceras	produced	0	0	1	0
producerar	producing	0	0	1	0
producerar	produces	0	0	1	0
köpa	purchase	0	0	1	1
köpa	buy	0	0	1	1
köpa	purchasing	0	0	1	0
grekisk	greek	0	0	1	1
producerat	produced	0	0	1	0
introducerade	introduced	0	0	1	0
producerade	produced	0	0	1	0
olycka	incident	0	0	1	0
olycka	accident	0	0	1	1
olycka	disaster	0	0	1	1
tro	believing	0	0	1	0
tro	think	0	0	1	1
budskap	message	0	0	1	1
graviditet	pregnancy	0	0	1	1
erkänt	recognized	0	0	1	0
blodet	the blood	0	0	1	0
blodet	blood	0	0	1	0
denne	his	0	0	1	0
denne	that he	0	0	1	0
denne	he	0	0	1	1
denna	that	0	0	1	0
uppehåll	residence	0	0	1	0
uppehåll	pause	0	0	1	1
uppehåll	hiatus	0	0	1	0
några	few	0	0	1	0
några	a few	0	0	1	0
enstaka	occasional	0	0	1	1
enstaka	single	0	0	1	1
england	england	0	0	1	1
bestämt	decided	0	0	1	1
bestämt	particularly	0	0	1	0
bestäms	determined	0	0	1	0
bestäms	is decided	0	0	1	0
slutgiltiga	final	0	0	1	0
doser	dose	0	0	1	0
operation	operation	0	0	1	1
återta	retake	0	0	1	0
återta	regain	0	0	1	0
återta	reclaim	0	0	1	0
finner	found	0	0	1	0
finner	finds	0	0	1	0
förutsättning	provided	0	0	1	0
förutsättning	quantity provided	0	0	1	0
förutsättning	prerequisite	0	0	1	0
jul	christmas	0	0	1	1
kopplad	connected to	0	0	1	0
kopplad	connected	0	0	1	0
garvey	garvey	0	0	1	0
avgick	resigned	0	0	1	0
avgick	retired	0	0	1	0
research	research	0	0	1	0
norska	norwegian	0	0	1	0
sammanfattning	summary	0	0	1	1
kopplat	coupled; connected	0	0	1	0
kopplat	connected	0	0	1	0
kopplat	coupled	0	0	1	0
kopplas	connected	0	0	1	0
kopplas	coupled	0	0	1	0
highway	highway	0	0	1	0
medel	middle	0	0	1	0
medel	medium	0	0	1	0
sparken	park	0	0	1	0
sparken	gets fired	0	0	1	0
sparken	fired	0	0	1	0
alltmer	increasingly	0	0	1	1
alltmer	more and more	0	0	1	1
poeter	poets	0	0	1	0
driver	run	0	0	1	0
driver	driver	0	0	1	1
driver	drive	0	0	1	0
kostade	cost	0	0	1	0
röra	move	0	0	1	1
poeten	poet	0	0	1	0
poeten	the poet	0	0	1	0
teknologi	technology	0	0	1	1
definition	defined	0	0	1	0
definition	definition	0	0	1	1
påverkad	affected	0	0	1	1
påverkad	influence	0	0	1	0
påverkad	influenced	0	0	1	0
kategorikrigsåret	category war years	0	0	1	0
gatorna	the streets	0	0	1	0
gatorna	streets	0	0	1	0
påverkan	impact	0	0	1	1
påverkan	influence	0	0	1	1
påverkar	affecting	0	0	1	0
påverkas	affected	0	0	1	0
påverkat	influenced	0	0	1	0
påverkat	affected	0	0	1	0
w	w	0	0	1	0
ägande	ownership	0	0	1	0
ägande	owning	0	0	1	1
föräldrar	parents	0	0	1	1
innebörd	meaning	0	0	1	0
innebörd	in meaning	0	0	1	0
vägarna	paths	0	0	1	0
vägarna	roads (roadways)	0	0	1	0
principen	the principal	0	0	1	0
principen	principle	0	0	1	0
bidragit	contributed	0	0	1	0
number	number	0	0	1	0
foten	foot	0	0	1	0
skiftande	shifting	0	0	1	1
spekulationer	speculation	0	0	1	0
spekulationer	speculations	0	0	1	0
gemensamma	joint	0	0	1	0
gemensamma	common	0	0	1	0
avel	breeding	0	0	1	1
avel	breed	0	0	1	0
liknas	compared to	0	0	1	0
liknas	likened	0	0	1	0
liknar	similar	0	0	1	0
liknar	similar to those	0	0	1	0
tove	tove	0	0	1	0
utökade	expanded	0	0	1	0
utökade	increased	0	0	1	0
saint	saint	0	0	1	0
natur	nature	0	0	1	1
missade	failed	0	0	1	0
anställd	employed	0	0	1	0
anställd	hired	0	0	1	0
följer	resulting	0	0	1	0
tappade	lost	0	0	1	0
zeus	zeus	0	0	1	1
striderna	the battles	0	0	1	0
striderna	fighting	0	0	1	0
förvaltning	management	0	0	1	1
förvaltning	administration	0	0	1	1
zeppelin	zeppelin	0	0	1	0
moder	parent	0	0	1	1
moder	mother	0	0	1	1
bidrog	contribute	0	0	1	0
bidrog	contributed	0	0	1	0
obama	obama	0	0	1	0
organiseras	organizes	0	0	1	0
organiseras	organized	0	0	1	0
organiserat	structured	0	0	1	0
niklas	niklas	0	0	1	0
koncentrerade	concentrated	0	0	1	0
koncentrerade	koncentrerade	0	0	1	0
marknadsekonomi	market economy	0	0	1	0
marknadsekonomi	market	0	0	1	0
freud	freud	0	0	1	0
organiserad	organised	0	0	1	0
organiserad	organized	0	0	1	1
hyde	hyde	0	0	1	0
rättigheter	rights	0	0	1	0
nikolaj	nikolaj	0	0	1	0
nikolaj	nicholas	0	0	1	0
inkluderas	include	0	0	1	0
inkluderas	is included	0	0	1	0
inkluderar	include	0	0	1	0
inkluderar	includes	0	0	1	0
möjligt	possible	0	0	1	0
generationen	generation	0	0	1	0
generationen	the generation	0	0	1	0
önskade	desired	0	0	1	0
önskade	wished	0	0	1	0
inkluderat	included	0	0	1	0
inkluderat	including	0	0	1	0
generationer	generation	0	0	1	0
generationer	generations	0	0	1	0
victoriasjön	victoria lake	0	0	1	0
victoriasjön	lake victoria	0	0	1	0
möjliga	possible	0	0	1	0
astronomin	the astronomy	0	0	1	0
astronomin	astronomy	0	0	1	0
förklaras	explained	0	0	1	0
förklarat	explained	0	0	1	0
förklarat	declare	0	0	1	0
visats	shown	0	0	1	0
visats	demonstrated	0	0	1	0
täcks	covered	0	0	1	0
täcks	covers	0	0	1	0
varianten	version	0	0	1	0
varianten	variant	0	0	1	0
norstedts	norstedt's	0	0	1	0
norstedts	norstedts	0	0	1	0
norstedts	collins	0	0	1	0
täckt	covered	0	0	1	1
täckt	coated	0	0	1	0
åtskilliga	several	0	0	1	1
kongokinshasa	kong kinshasa	0	0	1	0
kongokinshasa	democratic republic of the congo	0	0	1	0
kongokinshasa	congo kinshasa	0	0	1	0
fördraget	the treaty	0	0	1	0
fördraget	treaty	0	0	1	0
varianter	variants	0	0	1	0
varianter	varieties	0	0	1	0
varianter	diversities	0	0	1	0
täcka	cover	0	0	1	1
täcka	thank	0	0	1	0
vinterspelen	winter games	0	0	1	0
arabisk	arabic	0	0	1	1
försöka	try	0	0	1	1
försöka	attempt	0	0	1	1
sydostasien	south east asia	0	0	1	0
sydostasien	southeast asia	0	0	1	0
brooklyn	brooklyn	0	0	1	0
männen	the men	0	0	1	0
männen	men	0	0	1	0
plan	flat	0	0	1	1
plan	level	0	0	1	1
missnöje	miss our pleasure	0	0	1	0
missnöje	dissatisfaction	0	0	1	1
kombinationer	combinations	0	0	1	0
arter	species	0	0	1	0
utsattes	subjected	0	0	1	0
utsattes	were exposed	0	0	1	0
utsattes	exposed	0	0	1	0
cover	cover	0	0	1	0
kanalen	the channel	0	0	1	0
kanalen	channel	0	0	1	0
kanaler	channels	0	0	1	0
arten	species	0	0	1	0
kombinationen	the combination	0	0	1	0
kombinationen	combination	0	0	1	0
källan	source	0	0	1	0
källan	kallan	0	0	1	0
källan	the source	0	0	1	0
golf	golf	0	0	1	1
häst	horse	0	0	1	1
häst	haste	0	0	1	0
häst	equine	0	0	1	0
gold	gold	0	0	1	0
fackföreningar	unions	0	0	1	0
omfattade	included	0	0	1	0
omfattade	covered	0	0	1	0
berömd	famous	0	0	1	1
våld	violence	0	0	1	1
våld	force	0	0	1	1
presidentens	the president's	0	0	1	0
presidentens	president	0	0	1	0
presidentens	the presidents	0	0	1	0
uppförande	construction	0	0	1	1
uppförande	code	0	0	1	0
uppförande	behavior	0	0	1	1
detalj	detail	0	0	1	1
praktiken	effectively	0	0	1	0
praktiken	practice	0	0	1	0
praktiken	practically	0	0	1	0
berömt	famous	0	0	1	0
berömt	praised	0	0	1	0
falskt	false	0	0	1	0
existensen	existence	0	0	1	0
betydelser	meanings	0	0	1	0
betydelser	values	0	0	1	0
observatörer	observers	0	0	1	0
wayne	wayne	0	0	1	0
betydelsen	the meaning	0	0	1	0
betydelsen	significance	0	0	1	0
kontor	office	0	0	1	1
karakteristiska	characteristic	0	0	1	0
européer	europeans	0	0	1	0
genomgick	underwent	0	0	1	0
gratis	free	0	0	1	1
evolutionen	evolution	0	0	1	0
evolutionen	the evolution	0	0	1	0
tekniken	techinque	0	0	1	0
tekniken	art	0	0	1	0
tekniken	the technology	0	0	1	0
tekniker	technician	0	0	1	1
stätta	stood	1	0	1	0
stätta	created	1	0	1	0
stätta	ladder	1	1	0	0
stätta	stiles	1	1	0	0
stätta	start	1	0	1	0
stätta	stile	1	1	0	1
stätta	allow	1	0	1	0
stätta	tile	1	1	0	0
utbildningen	education	0	0	1	0
återvänt	atervant	0	0	1	0
återvänt	returned	0	0	1	0
återvänt	returning	0	0	1	0
crüe	crüe	0	0	1	0
tanken	the thought	0	0	1	0
tanken	idea	0	0	1	0
ledare	conductors	0	0	1	0
ledare	leader	0	0	1	1
bytet	the exchange	0	0	1	0
bytet	change	0	0	1	0
byter	changing	0	0	1	0
byter	changes	0	0	1	0
byter	exchanges	0	0	1	0
rösten	voice	0	0	1	0
rösten	the voice	0	0	1	0
rösten	rust	0	0	1	0
byten	byte	0	0	1	0
fotbeklädnad	chaussure	1	0	1	0
fotbeklädnad	foot gear	1	0	1	0
fotbeklädnad	chausurre	1	0	1	0
fotbeklädnad	shoewear	1	0	1	0
fotbeklädnad	footwear	1	1	0	1
fotbeklädnad	replacement	1	0	1	0
river	tear	0	0	1	0
river	river	0	0	1	0
avled	died	0	0	1	0
avled	deceased	0	0	1	0
nietzsches	nietzsche	0	0	1	0
nietzsches	nietzsche's	0	0	1	0
hällristning	halristning	1	0	1	0
hällristning	petroglyph	1	1	0	1
hällristning	rock	1	0	1	0
hällristning	stone carving	1	0	1	0
hällristning	agency	1	0	1	0
hällristning	rock engraving	1	0	1	0
hällristning	chives	1	0	1	0
hällristning	rock carvings	1	1	0	0
hällristning	n/a	1	0	1	0
hällristning	agencies	1	0	1	0
hällristning	rock carving	1	1	0	0
hällristning	rock engravings	1	0	1	0
hällristning	venom snooping	1	0	1	0
ser	see	0	0	1	0
ser	sees	0	0	1	0
koranen	the koran	0	0	1	0
koranen	the quran	0	0	1	0
sex	six	0	0	1	1
sed	sed	0	0	1	0
sed	thirst	0	0	1	0
psykologiska	psychological	0	0	1	0
uppkomsten	onset	0	0	1	0
uppkomsten	origin	0	0	1	0
sen	then	0	0	1	1
sen	since	0	0	1	1
sorters	kinds	0	0	1	0
sorters	kinds of	0	0	1	0
institutet	institute	0	0	1	0
institutet	the institution	0	0	1	0
project	project	0	0	1	0
äktenskap	the marriage	0	0	1	0
äktenskap	marriage	0	0	1	1
guinea	guinea	0	0	1	1
neutralitet	neutrality	0	0	1	1
neutralitet	neutral	0	0	1	0
antarktis	antarctica	0	0	1	1
antarktis	antarctic	0	0	1	1
fission	fission	0	0	1	1
sändebud	envoy	0	0	1	1
sändebud	messenger	0	0	1	0
alqaida	al-qaida	0	0	1	0
alqaida	al-qaeda	0	0	1	0
rita	paint	0	0	1	0
rita	draw	0	0	1	1
rita	drawing	0	0	1	0
europe	europe	0	0	1	0
europa	europe	0	0	1	1
europa	european	0	0	1	0
medveten	aware	0	0	1	1
medveten	conscious	0	0	1	1
avvikelser	abnormalities	0	0	1	0
avvikelser	deviations	0	0	1	0
avvikelser	derivations	0	0	1	0
medvetet	consciously	0	0	1	1
medvetet	conscious	0	0	1	0
näringslivet	economic life	0	0	1	0
näringslivet	industrial life	0	0	1	0
näringslivet	business	0	0	1	0
tävlingen	competition	0	0	1	0
tävlingen	contest	0	0	1	0
fame	fame	0	0	1	0
stadsdel	city district	0	0	1	0
stadsdel	neighborhood	0	0	1	0
stadsdel	district	0	0	1	1
utkom	issued	0	0	1	0
utkom	published	0	0	1	0
utkom	(was) issued	0	0	1	0
kategorimän	category: men	0	0	1	0
kategorimän	category men	0	0	1	0
släpptes	released	0	0	1	0
släpptes	was released	0	0	1	0
forskare	researcher	0	0	1	1
forskare	researchers	0	0	1	0
forskare	scientists	0	0	1	0
medicinering	medication	0	0	1	0
last	load	0	0	1	1
messias	messiah	0	0	1	1
dödsoffer	victim	0	0	1	1
dödsoffer	death victim	0	0	1	0
dödsoffer	casualty	0	0	1	0
halmstads	straw city	0	0	1	0
halmstads	halmstad's	0	0	1	0
kopia	copy	0	0	1	1
eftervärlden	posterity	0	0	1	0
eftervärlden	the world	0	0	1	0
kejsardömet	empire	0	0	1	0
samma	the same	0	0	1	1
samma	same	0	0	1	1
transeuropeiska	trans-european	0	0	1	0
transeuropeiska	transeuropean	0	0	1	0
bell	bell	0	0	1	0
olle	olle	0	0	1	0
långtgående	far-reaching	0	0	1	0
kriser	crises	0	0	1	0
church	church	0	0	1	0
allierade	allied	0	0	1	0
allierade	allies	0	0	1	0
språkets	the language's	0	0	1	0
språkets	language	0	0	1	0
föreningar	associations	0	0	1	0
föreningar	organizations	0	0	1	0
föreningar	compounds	0	0	1	0
populärmusik	popular music	0	0	1	0
populärmusik	pop music	0	0	1	0
fått	was given	0	0	1	0
fått	with	0	0	1	0
sommaren	summer	0	0	1	0
sommaren	the summer	0	0	1	0
koalition	coalition	0	0	1	1
potentiellt	potential	0	0	1	0
kyrilliska	cyrillic	0	0	1	0
blod	blood	0	0	1	1
gällande	current	0	0	1	1
gällande	regarding	0	0	1	0
uppträda	act	0	0	1	1
uppträda	appear	0	0	1	1
uppträda	occur	0	0	1	0
beskrevs	was described	0	0	1	0
beskrevs	described	0	0	1	0
nivån	level	0	0	1	0
fire	fire	0	0	1	0
stadskärnan	town/city	0	0	1	0
stadskärnan	city bear man	0	0	1	0
stadskärnan	center	0	0	1	0
fira	celebrate	0	0	1	1
fritz	fritz	0	0	1	0
avrättningen	execution	0	0	1	0
avrättningen	the execution	0	0	1	0
fritt	free	0	0	1	1
systematik	systematics	0	0	1	0
systematik	systematic	0	0	1	0
handling	action	0	0	1	1
handling	act	0	0	1	1
projekt	project	0	0	1	1
knä	knee	0	0	1	1
knä	knees	0	0	1	0
budget	budget	0	0	1	1
guldbollen	the ball	0	0	1	0
guldbollen	golden ball	0	0	1	0
guldbollen	guldbollen	0	0	1	0
robin	robin	0	0	1	0
pressen	press	0	0	1	0
pressen	the pres	0	0	1	0
real	real	0	0	1	1
österrikeungern	oster kingdom hungary	0	0	1	0
österrikeungern	austria-hungary	0	0	1	0
vägen	the road	0	0	1	0
vägen	road	0	0	1	0
arbete	work	0	0	1	1
arbete	work; labor	0	0	1	0
vol	v	0	0	1	0
målvakten	the goalkeeper	0	0	1	0
von	von	0	0	1	0
owen	owen	0	0	1	0
motors	engine's	0	0	1	0
motors	motor	0	0	1	0
titanic	titanic	0	0	1	0
lokaler	facilities	0	0	1	0
lokaler	studios	0	0	1	0
lokaler	place	0	0	1	0
väger	weighs	0	0	1	0
väger	weight	0	0	1	0
madagaskar	madagascar	0	0	1	1
utmärkande	characteristic	0	0	1	0
utmärkande	distinguishing	0	0	1	1
hovet	court	0	0	1	0
hovet	the court	0	0	1	0
kritiker	critics	0	0	1	0
kritiker	critiques	0	0	1	0
objekt	objects	0	0	1	1
objekt	object	0	0	1	1
närmade	approached	0	0	1	0
tecken	signs	0	0	1	0
tecken	characters	0	0	1	0
tecken	sign	0	0	1	1
barnet	child	0	0	1	0
omvandlar	converts	0	0	1	0
omvandlar	transmuted	0	0	1	0
skalet	shell	0	0	1	0
skalet	the shell	0	0	1	0
barnen	children	0	0	1	0
föreställningen	the idea	0	0	1	0
föreställningen	the concept	0	0	1	0
föreställningen	show	0	0	1	0
kritiken	criticism	0	0	1	0
kritiken	the criticism	0	0	1	0
kritiken	the critique	0	0	1	0
laddning	charge	0	0	1	1
kategoriavlidna	kategoriavlidna	0	0	1	0
kategoriavlidna	category deceased	0	0	1	0
debatter	debates	0	0	1	0
rådhus	townhouses	0	0	1	0
rådhus	town hall	0	0	1	1
rådhus	courthouse	0	0	1	0
republiken	the republic of	0	0	1	0
republiken	the republic	0	0	1	0
republiker	republics	0	0	1	0
grannlandet	neighboring	0	0	1	0
grannlandet	the neighbouring country	0	0	1	0
kring	on	0	0	1	0
kring	around	0	0	1	0
ledarskap	leadership	0	0	1	1
fyra	four	0	0	1	1
vargar	wolves	0	0	1	0
euro	euro	0	0	1	0
normala	normal	0	0	1	0
västtyskland	västttyskland	0	0	1	0
västtyskland	west germany	0	0	1	1
normalt	normally	0	0	1	1
normalt	normal	0	0	1	0
person	person	0	0	1	1
kelly	kelly	0	0	1	0
johan	john	0	0	1	0
johan	johan	0	0	1	0
kontakter	contact	0	0	1	0
kontakter	contacts	0	0	1	0
finansiellt	financial	0	0	1	0
konkret	specific	0	0	1	0
konkret	concrete	0	0	1	1
tunnelbana	subway	0	0	1	1
telegram	telegram	0	0	1	1
koprolali	coprolalia	1	1	0	0
koprolali	number	1	0	1	0
koprolali	coporolalia	1	0	1	0
stockholms	stockholm's	0	0	1	0
stockholms	stockholm	0	0	1	0
trädgård	garden	0	0	1	1
webbkällor	websources	0	0	1	0
webbkällor	webbkällor	0	0	1	0
webbkällor	web sources	0	0	1	0
finansiella	financial	0	0	1	0
kontakten	connector	0	0	1	0
kontakten	the contact	0	0	1	0
kontakten	conntact	0	0	1	0
mandat	mandate	0	0	1	1
fascistiska	fascist	0	0	1	0
fascistiska	fascistic	0	0	1	0
rebecca	rebecca	0	0	1	0
festivalen	festival	0	0	1	0
festivalen	the festival	0	0	1	0
återkommer	recurs	0	0	1	0
återkommer	will return	0	0	1	0
återkommer	returning	0	0	1	0
läge	mode	0	0	1	1
läge	location	0	0	1	1
symbolisk	nominal	0	0	1	1
symbolisk	symbolic	0	0	1	1
festivaler	festivals	0	0	1	0
läror	teachings	0	0	1	0
tomas	tomas	0	0	1	0
australia	australia	0	0	1	0
format	format	0	0	1	1
format	shaped	0	0	1	0
teologiska	theological	0	0	1	0
här	this; here	0	0	1	0
här	is	0	0	1	0
här	here	0	0	1	1
nämligen	namely	0	0	1	1
melker	melker	0	0	1	0
avvisar	reject	0	0	1	0
skara	city in south-central sweden (uppland)	0	0	1	0
skara	crowd	0	0	1	0
samarbete	collaboration	0	0	1	1
samarbete	co	0	0	1	0
ivar	ivar	0	0	1	0
samarbeta	collaborate	0	0	1	1
samarbeta	co	0	0	1	0
samarbeta	cooperate	0	0	1	1
upptäckter	discoveries	0	0	1	0
upptäckter	discovery	0	0	1	0
upptäcktes	discovered	0	0	1	0
upptäcktes	(was) discovered	0	0	1	0
funnit	found	0	0	1	0
skarp	sharp	0	0	1	1
skarp	crisp	0	0	1	0
informationen	the information	0	0	1	0
västeuropa	western europe	0	0	1	1
västeuropa	west europe	0	0	1	0
upptäckten	the discovery	0	0	1	0
upptäckten	discovery	0	0	1	0
patrick	patrick	0	0	1	0
ivan	ivan	0	0	1	0
alexandra	alexandra	0	0	1	0
evangelierna	gospels	0	0	1	0
evangelierna	the gospels	0	0	1	0
östersjön	baltic	0	0	1	0
östersjön	balticsea	0	0	1	0
vojvodina	voyvodina	0	0	1	0
vojvodina	vojvodina	0	0	1	0
lenin	lenin	0	0	1	0
långstrump	hose drumstick	0	0	1	0
långstrump	longstocking	0	0	1	0
rörelse	movement	0	0	1	1
saknar	lacks	0	0	1	0
saknar	lack(-s)	0	0	1	0
saknar	missing	0	0	1	0
saknas	missing	0	0	1	0
utvecklades	developed	0	0	1	0
utvecklades	(was) developed	0	0	1	0
påstådda	said	0	0	1	0
påstådda	alleged	0	0	1	0
avskaffade	abolished	0	0	1	0
avskaffade	absolished	0	0	1	0
wallenstein	wallenstein	0	0	1	0
köra	run	0	0	1	0
köra	drive	0	0	1	1
genomfördes	completed	0	0	1	0
genomfördes	was	0	0	1	0
genomfördes	was carried out	0	0	1	0
brasilianska	brasilian	0	0	1	0
brasilianska	brazilian	0	0	1	0
största	biggest	0	0	1	0
största	maximum	0	0	1	0
största	largest	0	0	1	0
trafiken	traffic	0	0	1	0
trafiken	the traffic	0	0	1	0
turnerade	toured	0	0	1	0
religion	religion	0	0	1	1
körs	driven	0	0	1	0
körs	running	0	0	1	0
körs	being driven	0	0	1	0
drogmissbruk	drug abuse	0	0	1	0
drogmissbruk	drug addiction	0	0	1	0
drogmissbruk	drug	0	0	1	0
drogmissbruk	substance abuse	0	0	1	0
vacker	beautiful	0	0	1	1
överst	top	0	0	1	0
överst	at the top; uppermost	0	0	1	0
nybildade	newly formed	0	0	1	0
nybildade	newly established	0	0	1	0
ugandas	of uganda	0	0	1	0
ugandas	uganda	0	0	1	0
bl	bl	0	0	1	0
bl	short of "bland" - in the context: bl. a (bland annat) = among others	0	0	1	0
ifråga	with regards to	0	0	1	0
ifråga	in question	0	0	1	0
ifråga	challenged	0	0	1	0
krita	chalk	0	0	1	1
bo	living	0	0	1	0
belägen	located	0	0	1	1
belägen	situated	0	0	1	1
belägen	disposed	0	0	1	0
bk	bk	0	0	1	0
plocka	pick	0	0	1	1
engelska	england	0	0	1	0
engelska	english	0	0	1	1
bokstav	character	0	0	1	1
bokstav	letter	0	0	1	1
ordning	system	0	0	1	0
bildat	formed	0	0	1	0
santa	santa	0	0	1	0
by	by	0	0	1	0
by	village	0	0	1	1
riksförbundet	national association	0	0	1	0
ideologin	ideology	0	0	1	0
ideologin	the ideology	0	0	1	0
återvänder	returns	0	0	1	0
återvänder	atervander	0	0	1	0
upprätta	establish	0	0	1	1
upprätta	up	0	0	1	0
dagligen	day	0	0	1	0
dagligen	daily	0	0	1	1
gemenskaperna	communities	0	0	1	0
gemenskaperna	community	0	0	1	0
aggressiv	aggressive	0	0	1	1
umgänge	company	0	0	1	1
umgänge	intercourse	0	0	1	1
stuart	stuart	0	0	1	0
fungerande	functioning	0	0	1	0
fungerande	working	0	0	1	0
fungerande	effective	0	0	1	0
papper	paper	0	0	1	1
texterna	text	0	0	1	0
inte	not	0	0	1	1
inta	taken	0	0	1	0
colorado	colorado	0	0	1	0
syret	the oxygen	0	0	1	0
syret	oxygen	0	0	1	0
tyvärr	unfortunately	0	0	1	1
hemingway	hemingway	0	0	1	0
kravet	requirement	0	0	1	0
kravet	the demand	0	0	1	0
spridas	spread	0	0	1	0
spridas	disseminated	0	0	1	0
kraven	the demands	0	0	1	0
kraven	requirements	0	0	1	0
uppkallad	named	0	0	1	0
seger	victory	0	0	1	1
jönsson	johnsson	0	0	1	0
jönsson	jönsson	0	0	1	0
veckor	weeks	0	0	1	0
kategorimusikgrupper	category of music groups	0	0	1	0
svårt	hard	0	0	1	0
svårt	black	0	0	1	0
svårt	difficult	0	0	1	0
inlägg	post	0	0	1	0
framträdde	appeared	0	0	1	0
framträdde	emerged	0	0	1	0
u+	u +	0	0	1	0
samerna	sami	0	0	1	0
samerna	the lapp	0	0	1	0
svåra	answering	0	0	1	0
svåra	difficult	0	0	1	0
knuten	tied to	0	0	1	0
knuten	bound	0	0	1	0
knuten	knot	0	0	1	0
fattigdom	poverty	0	0	1	1
fattigdom	fattidom	0	0	1	0
poster	positions	0	0	1	0
poster	post offices	0	0	1	0
rött	cane	0	0	1	0
rött	red	0	0	1	1
betyda	mean	0	0	1	1
begreppet	the term	0	0	1	0
begreppet	term	0	0	1	0
begreppet	concept	0	0	1	0
posten	post	0	0	1	0
posten	the position	0	0	1	0
atom	atomic	0	0	1	0
atom	atom	0	0	1	1
kritisk	critical	0	0	1	1
line	line	0	0	1	0
lovade	promised	0	0	1	0
heinrich	heinrich	0	0	1	0
röster	votes	0	0	1	0
katoliker	catholics	0	0	1	0
cia	cia	0	0	1	0
ut	out; up	0	0	1	0
ut	out	0	0	1	1
godkännande	approval	0	0	1	1
godkännande	authorization	0	0	1	0
eddie	eddie	0	0	1	0
us	oss	0	0	1	0
ur	from	0	0	1	1
ur	out	0	0	1	0
konventionella	conventional	0	0	1	0
distrikt	district	0	0	1	1
uk	uk	0	0	1	0
galaxer	galaxies	0	0	1	0
högkvarter	headquarters	0	0	1	1
högkvarter	head quarter	0	0	1	0
testamente	testament	0	0	1	1
testamente	will	0	0	1	1
testamente	wills	0	0	1	0
erics	erics	0	0	1	0
lägst	lowest	0	0	1	1
lägst	lowermost	0	0	1	1
pernilla	pernilla	0	0	1	0
diverse	some	0	0	1	0
diverse	miscellaneous	0	0	1	1
utbyggt	develpoed	0	0	1	0
utbyggt	built	0	0	1	0
utbyggt	extended	0	0	1	0
makedonska	macedonian	0	0	1	0
makedonska	makedonish	0	0	1	0
nationalism	nationalism	0	0	1	1
inblandning	incorporation	0	0	1	0
inblandning	involvement	0	0	1	1
väder	weather	0	0	1	1
matematiken	mathematics	0	0	1	0
gestalter	beings	0	0	1	0
gestalter	figures	0	0	1	0
ingått	been part of	0	0	1	0
ingått	entered	0	0	1	0
ingått	entered into	0	0	1	0
skrivits	down	0	0	1	0
skrivits	srivits	0	0	1	0
skrivits	been written	0	0	1	0
nordafrika	north africa	0	0	1	0
matematiker	mathematician	0	0	1	1
existerade	existed	0	0	1	0
existerade	existing	0	0	1	0
upplaga	edition	0	0	1	1
upplaga	uppalaga	0	0	1	0
upplaga	submission	0	0	1	0
individuella	individual	0	0	1	0
besegra	defeat	0	0	1	1
dominerades	was dominated	0	0	1	0
dominerades	dominated	0	0	1	0
radikala	radical	0	0	1	0
lucia	lucia	0	0	1	0
konstantinopel	constantinople	0	0	1	0
riskerar	could	0	0	1	0
riskerar	risks	0	0	1	0
riskerar	there is a risk	0	0	1	0
nästan	almost	0	0	1	1
nästan	close	0	0	1	0
springsteen	springsteen	0	0	1	0
radikalt	radical	0	0	1	0
radikalt	radically	0	0	1	1
hells	hells	0	0	1	0
land	country	0	0	1	1
passagerarna	passengers	0	0	1	0
passagerarna	the passengers	0	0	1	0
målade	painted	0	0	1	0
symtom	symptoms	0	0	1	0
symtom	symptom	0	0	1	0
produkt	product	0	0	1	1
texten	text	0	0	1	0
texten	the text	0	0	1	0
sawyer	sawyer	0	0	1	0
texter	texts	0	0	1	0
båtar	boats	0	0	1	0
majs	corn	0	0	1	1
persbrandt	persbrandt	0	0	1	0
koloniserades	is colonized	0	0	1	0
koloniserades	colonized	0	0	1	0
störtades	overthrew	0	0	1	0
störtades	overthrown	0	0	1	0
störtades	was overthrown	0	0	1	0
utökat	extended	0	0	1	0
utökat	expanded	0	0	1	0
anorektiker	anorectics	0	0	1	0
anorektiker	anorexic	0	0	1	0
anorektiker	anorectic	0	0	1	0
turkisk	turkish	0	0	1	1
dyraste	most expensive	0	0	1	0
sena	late	0	0	1	0
young	small	0	0	1	0
listade	listed	0	0	1	0
sydväst	southwest	0	0	1	1
dickinson	dickinson	0	0	1	0
monoteistiska	monotheistic	0	0	1	0
sent	late	0	0	1	1
garden	garden	0	0	1	0
dagsläget	present situation	0	0	1	0
dagsläget	current situation	0	0	1	0
någorlunda	fairly	0	0	1	1
någorlunda	somewhat	0	0	1	0
hustru	wife	0	0	1	1
palestinier	palestinians	0	0	1	0
palestinier	palestinian	0	0	1	1
kommunistiska	communistic	0	0	1	0
kommunistiska	communist	0	0	1	0
drogen	the drug	0	0	1	0
drogen	drug	0	0	1	0
vinner	gaining	0	0	1	0
vinner	wins	0	0	1	0
vinner	win	0	0	1	0
magic	magic	0	0	1	0
dök	appeared	0	0	1	0
dök	turned	0	0	1	0
dök	dove	0	0	1	0
omvänt	reversed	0	0	1	0
omvänt	vice versa	0	0	1	1
harbor	harbor	0	0	1	0
eva	eva	0	0	1	0
tre	three	0	0	1	1
jobbet	work	0	0	1	0
jobbet	the job	0	0	1	0
därvid	thus; thusly; then	0	0	1	0
därvid	therewith	0	0	1	0
därvid	in so doing	0	0	1	0
romerska	roman	0	0	1	0
romerske	roman	0	0	1	0
död	death	0	0	1	1
död	dod	0	0	1	0
död	dead	0	0	1	1
erkänd	acknowledged	0	0	1	1
erkänd	recognized	0	0	1	1
opinionen	opinion	0	0	1	0
leonardo	leonardo	0	0	1	0
bolsjevikerna	bolsevikema	0	0	1	0
bolsjevikerna	bolsheviks	0	0	1	0
bolsjevikerna	the bolsheviks	0	0	1	0
nordvästra	northwest	0	0	1	0
nordvästra	north western	0	0	1	0
regelbundna	regular	0	0	1	0
video	video	0	0	1	1
dessförinnan	before (that)	0	0	1	0
dessförinnan	before	0	0	1	0
victor	victor	0	0	1	0
antog	adopted	0	0	1	0
index	index	0	0	1	1
högskolan	hogs school	0	0	1	0
högskolan	university	0	0	1	0
högskolan	college	0	0	1	0
nevada	nevada	0	0	1	0
expressen	expressen	0	0	1	0
anton	anton	0	0	1	0
byrå	bureau	1	1	0	1
fritid	free time	1	1	0	0
fritid	record	1	0	1	0
fritid	recreational	1	0	1	0
fritid	leisure	1	1	0	1
fritid	records	1	0	1	0
fritid	leisure time	1	1	0	1
fritid	freetime	1	1	0	0
fritid	spare time	1	0	1	1
fritid	leisure time; spare time	1	0	1	0
indiens	india's	0	0	1	0
indiens	indias	0	0	1	0
richmond	richmond	0	0	1	0
birk	brik	0	0	1	0
birk	birk	0	0	1	0
indian	indian	0	0	1	1
ledande	conductive	0	0	1	1
ledande	leading	0	0	1	1
läkare	doctor	0	0	1	1
läkare	doctors	0	0	1	0
försökt	tried	0	0	1	0
mästare	master	0	0	1	1
mästare	champion	0	0	1	1
led	step	0	0	1	0
led	suffered	0	0	1	0
lee	lee	0	0	1	0
lyckades	managed	0	0	1	0
lyckades	succeeded	0	0	1	0
leo	leo	0	0	1	0
les	les	0	0	1	0
let	cleanly	0	0	1	0
lev	live	0	0	1	0
lev	lev	0	0	1	0
talang	talent	0	0	1	1
begravd	buried	0	0	1	1
tegel	brick	0	0	1	1
casino	casino	0	0	1	0
försörjning	sustention	0	0	1	0
försörjning	sustentation	0	0	1	0
försörjning	supply	0	0	1	0
trä	tra	0	0	1	0
trä	wood	0	0	1	1
fängelsestraff	imprisonment	0	0	1	1
fängelsestraff	prison	0	0	1	0
förlust	loss	0	0	1	1
tillkom	hold back	0	0	1	0
tillkom	resided	0	0	1	0
insulin	insulin	0	0	1	1
opinion	opinion	0	0	1	0
dör	dies	0	0	1	0
dör	die	0	0	1	0
dålig	poor	0	0	1	1
artisterna	aristerna	0	0	1	0
artisterna	artists	0	0	1	0
emot	vis	0	0	1	0
emot	against	0	0	1	1
åker	go	0	0	1	0
åker	treats	0	0	1	0
åker	field; going	0	0	1	0
oxenstierna	the oxenstierna	0	0	1	0
oxenstierna	oxenstierna	0	0	1	0
mening	meaning	0	0	1	1
mening	meanings	0	0	1	0
mening	sentence	0	0	1	1
fotosyntesen	photosynthesis	0	0	1	0
anatolien	anatolia	0	0	1	0
tillägg	addition	0	0	1	1
tillägg	appendix	0	0	1	0
känd	known	0	0	1	1
känd	unknown	0	0	1	0
känd	famous	0	0	1	1
varmare	heater	0	0	1	0
varmare	warmer	0	0	1	0
illegal	illicit	0	0	1	1
illegal	illegal	0	0	1	1
överföra	transmit	0	0	1	1
överföra	transfer	0	0	1	1
hemlig	secret	0	0	1	1
elever	students	0	0	1	0
rätt	steering wheel	0	0	1	0
rätt	right	0	0	1	1
rätt	entitled	0	0	1	0
fjärde	fourth	0	0	1	1
känt	known	0	0	1	0
känt	famous	0	0	1	0
känt	side	0	0	1	0
klaviatur	keyboard	0	0	1	1
förändringen	the change	0	0	1	0
förändringen	change	0	0	1	0
förändringen	change.	0	0	1	0
överförs	is transferred	0	0	1	0
överförs	transfered	0	0	1	0
fält	field	0	0	1	1
orkester	orchestra	0	0	1	1
tillkännagav	announced	0	0	1	0
föredrog	prefered	0	0	1	0
föredrog	preferred	0	0	1	0
projektet	project	0	0	1	0
träffas	meet	0	0	1	1
träffas	reached	0	0	1	0
herbert	herbert	0	0	1	0
siffror	figures	0	0	1	0
siffror	numbers	0	0	1	0
samspel	interaction	0	0	1	0
samspel	teamwork	0	0	1	1
ytterst	very; extremely	0	0	1	0
ytterst	highly	0	0	1	0
villor	houses	0	0	1	0
villor	villas	0	0	1	0
edwall	edwall	0	0	1	0
lokalt	locally	0	0	1	0
lokalt	local	0	0	1	0
bidraget	contribution	0	0	1	0
bidraget	grant	0	0	1	0
benämns	designated	0	0	1	0
benämns	is mentioned	0	0	1	0
advokat	bar	0	0	1	0
advokat	lawyer	0	0	1	1
ortodoxa	orthodox	0	0	1	0
lokala	local	0	0	1	0
befolkningstillväxten	population growth	0	0	1	0
befolkningstillväxten	the growth of population	0	0	1	0
befolkningstillväxten	the population growth	0	0	1	0
giftermål	marriage	0	0	1	1
giftermål	marrige	0	0	1	0
peka	point (at; to; in)	0	0	1	0
peka	point	0	0	1	1
höll	held	0	0	1	0
höll	hold	0	0	1	0
höll	gave	0	0	1	0
frånvaro	absent	0	0	1	0
frånvaro	absence	0	0	1	1
sekel	centuries	0	0	1	0
sekel	century	0	0	1	1
process	process	0	0	1	1
artiklar	items	0	0	1	0
etta	number one	0	0	1	0
etta	one	0	0	1	1
etta	first	0	0	1	0
tryckta	printed	0	0	1	0
high	high	0	0	1	0
översätts	translated	0	0	1	0
översätts	translate	0	0	1	0
översätts	is translated	0	0	1	0
syre	oxygen	0	0	1	1
hercegovina	herzegovina	0	0	1	0
från	from	0	0	1	1
halmstad	halmstad	0	0	1	0
halmstad	halmstad's	0	0	1	0
gitarr	guitar	0	0	1	1
gitarr	guitarr	0	0	1	0
anländer	arrive	0	0	1	0
anländer	arrives	0	0	1	0
delad	shared	0	0	1	1
delad	divided	0	0	1	1
militärer	military	0	0	1	0
militärer	soldiers	0	0	1	0
latinska	latin	0	0	1	0
militären	military	0	0	1	0
militären	the military	0	0	1	0
hormoner	hormons	0	0	1	0
hormoner	hormones	0	0	1	0
överens	in agreement	0	0	1	0
överens	agree	0	0	1	0
delas	shared	0	0	1	0
delas	divided	0	0	1	0
delar	proportions	0	0	1	0
delar	parts	0	0	1	0
delat	shared	0	0	1	0
delat	divided	0	0	1	0
besläktat	related to	0	0	1	0
besläktat	related	0	0	1	0
bränder	fires	0	0	1	0
brändes	burned	0	0	1	0
brändes	burnt	0	0	1	0
gunwer	gunwer	0	0	1	0
amerika	american	0	0	1	0
amerika	america	0	0	1	1
djurens	the animals	0	0	1	0
djurens	animal	0	0	1	0
profeten	prophet	0	0	1	0
profeten	the prophet	0	0	1	0
insatser	action	0	0	1	0
regeringsmakten	govermental power	0	0	1	0
regeringsmakten	government power	0	0	1	0
bål	prom	0	0	1	0
bål	torso	0	0	1	1
förbättrade	improved	0	0	1	0
förbättrade	improve	0	0	1	0
slutsatser	conclusions	0	0	1	0
element	elements	0	0	1	0
lundgren	lundgren	0	0	1	0
nancy	nancy	0	0	1	0
kvinnliga	female	0	0	1	0
förblir	remains	0	0	1	0
förblir	remain	0	0	1	0
tätort	urban	0	0	1	0
tätort	conurbation	0	0	1	0
saknade	lacked	0	0	1	0
saknade	missed	0	0	1	0
saknade	missing	0	0	1	0
handboll	handball	0	0	1	1
diskar	disks	0	0	1	0
houston	houston	0	0	1	0
universiteten	universities	0	0	1	0
universiteten	the universities	0	0	1	0
bedöms	expected	0	0	1	0
bedöms	judged	0	0	1	0
bedöms	evaluated	0	0	1	0
hunnit	reached	0	0	1	0
hunnit	had	0	0	1	0
hunnit	had time to	0	0	1	0
universitetet	the university	0	0	1	0
universitetet	university	0	0	1	0
bedöma	judge; decide	0	0	1	0
bedöma	assessment	0	0	1	0
solvinden	the solar wind	0	0	1	0
solvinden	solar wind	0	0	1	0
eliten	the elite	0	0	1	0
eliten	elite	0	0	1	0
uppdelat	divided	0	0	1	0
uppdelat	split	0	0	1	0
möjligen	possibly	0	0	1	1
möjligen	it may have	0	0	1	0
tecknet	the sign	0	0	1	0
tecknet	sign	0	0	1	0
uppdelad	divided	0	0	1	0
uppdelad	split	0	0	1	0
puerto	puerto	0	0	1	0
puerto	port	0	0	1	0
utifrån	from the outside	0	0	1	1
utifrån	from	0	0	1	0
ovanlig	unusual	0	0	1	1
ovanlig	rare	0	0	1	1
ovanlig	uncommon	0	0	1	1
konkurs	bankrupcy	0	0	1	0
konkurs	bankruptcy	0	0	1	1
bekant	known	0	0	1	1
bekant	acquaintance	0	0	1	0
böckerna	books	0	0	1	0
bryter	breaks	0	0	1	0
bryter	breaking; violating	0	0	1	0
österut	eastwards	0	0	1	1
österut	east	0	0	1	1
beståndsdelar	constituents	0	0	1	0
beståndsdelar	elements	0	0	1	0
ställa	make	0	0	1	0
ställa	set	0	0	1	1
ställa	installation	0	0	1	0
hemmaplan	home	0	0	1	0
hemmaplan	home turf; domestic (level)	0	0	1	0
dock	nevertheless	0	0	1	1
dock	however	0	0	1	1
kiss	kiss	0	0	1	0
kiss	view	0	0	1	0
indikerar	indicates	0	0	1	0
rotation	rotation	0	0	1	1
ställt	put	0	0	1	0
ställt	taken	0	0	1	0
ställt	set	0	0	1	0
ställs	is	0	0	1	0
ställs	stalls	0	0	1	0
huvuddelen	bulk	0	0	1	0
huvuddelen	main part	0	0	1	0
framföra	express	0	0	1	0
framföra	convey	0	0	1	1
symboliserar	symbolized	0	0	1	0
symboliserar	symbolizes	0	0	1	0
peking	beijing	0	0	1	0
peking	peking	0	0	1	1
bipolära	bipolar	0	0	1	0
benämning	term	0	0	1	1
benämning	name	0	0	1	1
benämning	title	0	0	1	0
kriminella	criminal	0	0	1	0
intressen	interests	0	0	1	1
smallwood	small wood	0	0	1	0
smallwood	smallwood	0	0	1	0
svårare	answering machine	0	0	1	0
svårare	harder	0	0	1	0
svårare	difficult	0	0	1	0
society	society	0	0	1	0
books	books	0	0	1	0
fjärdedel	quarter	0	0	1	1
fjärdedel	fourth	0	0	1	1
intresset	interests	0	0	1	0
intresset	the interest	0	0	1	0
intresset	interest	0	0	1	0
frac	fraction	0	0	1	0
konsubstantiation	no idea what it means	1	0	1	0
konsubstantiation	konsubstantiaion	1	0	1	0
konsubstantiation	korea	1	0	1	0
konsubstantiation	consubstantion	1	0	1	0
konsubstantiation	konsubstantiation	1	0	1	0
konsubstantiation	consubstantiation	1	1	0	0
konsubstantiation	con-substantiation	1	0	1	0
etymologi	etymology	0	0	1	1
matrix	matrix	0	0	1	0
borderline	borderline	0	0	1	0
billiga	cheap	0	0	1	0
utbildad	formed	0	0	1	0
utbildad	educated	0	0	1	0
enskilda	individual	0	0	1	0
anledningen	reason	0	0	1	0
anledningen	therefore	0	0	1	0
kapitalismens	capitalism	0	0	1	0
kapitalismens	capitalism's	0	0	1	0
marxistiska	marxist	0	0	1	0
undertecknades	signed	0	0	1	0
medföra	bring	0	0	1	1
medföra	imply; entail	0	0	1	0
medföra	result	0	0	1	0
medföra	lead; result in	0	0	1	0
redskap	device	0	0	1	0
redskap	tool	0	0	1	1
egenskaperna	the qualities	0	0	1	0
egenskaperna	properties	0	0	1	0
release	release	0	0	1	0
underverk	wonder	0	0	1	1
underverk	wonders	0	0	1	0
uppe	(on) top	0	0	1	0
uppe	top	0	0	1	0
uppe	up	0	0	1	1
uppe	above	0	0	1	0
lundin	lundin	0	0	1	0
återförening	reunion	0	0	1	1
själ	shawl	0	0	1	0
själ	soul	0	0	1	1
dubbel	double	0	0	1	1
önskan	desired	0	0	1	0
önskan	our dreams	0	0	1	0
david	david	0	0	1	0
blanda	mix	0	0	1	1
profeter	prophets	0	0	1	0
profeter	profets	0	0	1	0
önskar	desired	0	0	1	0
önskar	desiring to	0	0	1	0
önskar	wish	0	0	1	0
krets	sphere	0	0	1	1
krets	circuit	0	0	1	1
helst	rather	0	0	1	0
helst	anyone	0	0	1	0
helst	any time	0	0	1	0
förstärka	strengthen	0	0	1	1
förstärka	enhance	0	0	1	0
förnuftet	reason	0	0	1	0
förnuftet	the common sense	0	0	1	0
hussein	hussein	0	0	1	0
skillnad	difference	0	0	1	1
skillnad	unlike	0	0	1	0
sjukvård	health care	0	0	1	0
sjukvård	care	0	0	1	0
sjukvård	healthcare	0	0	1	0
playstation	playstation	0	0	1	0
komplicerade	konplicerade	0	0	1	0
komplicerade	complex	0	0	1	0
jesus	jesus	0	0	1	1
fågelhundar	bird dogs	0	0	1	0
muhammad	muhammad	0	0	1	0
sköttes	operated	0	0	1	0
sköttes	handled	0	0	1	0
nordkoreanska	north korean	0	0	1	0
studerade	studied	0	0	1	0
nationalistiska	nationalist	0	0	1	0
nationalistiska	nationalistic	0	0	1	0
förkortas	shortened	0	0	1	0
förkortas	abbreviated	0	0	1	0
förkortas	reduced	0	0	1	0
förkortat	shortened	0	0	1	0
förkortat	abbreviated	0	0	1	0
start	start	0	0	1	1
festival	festival	0	0	1	1
system	system	0	0	1	1
bygget	the construction	0	0	1	0
bygget	construction	0	0	1	0
syster	sister	0	0	1	1
hebreiska	hebrew	0	0	1	1
teatern	the theater	0	0	1	0
teatern	theater	0	0	1	0
blivit	become	0	0	1	0
blivit	was	0	0	1	0
osäkra	insecure	0	0	1	0
osäkra	uncertain	0	0	1	0
osäkra	doubtful	0	0	1	0
utbyggnad	development	0	0	1	1
utbyggnad	addition	0	0	1	0
utbyggnad	expansion	0	0	1	0
havet	sea	0	0	1	0
sömn	sleep	0	0	1	1
pristagare	laureate	0	0	1	0
pristagare	prizewinner	0	0	1	0
konservativ	conservative	0	0	1	1
haven	the seas	0	0	1	0
visdom	wisdom	0	0	1	1
hampa	hemp	0	0	1	1
samverkar	co-operating	0	0	1	0
samverkar	co	0	0	1	0
samverkar	co-operates	0	0	1	0
roberto	roberto	0	0	1	0
grundarna	founders	0	0	1	0
aktörer	players	0	0	1	0
aktörer	actors	0	0	1	0
roberts	roberts	0	0	1	0
låtit	let	0	0	1	0
låtit	ordered	0	0	1	0
låtit	had	0	0	1	0
reagans	reagan's	0	0	1	0
reagans	reagan	0	0	1	0
troende	believers	0	0	1	1
troende	faithful	0	0	1	0
vecka	week	0	0	1	1
jonatan	jonatan	0	0	1	0
jonatan	jonathan	0	0	1	0
dräkt	costume	0	0	1	1
dräkt	outfit	0	0	1	0
inre	inner	0	0	1	1
årsdag	anniversary	0	0	1	1
talrika	numerous	0	0	1	0
mänskligheten	humanity	0	0	1	1
mänskligheten	manskligheten	0	0	1	0
flygplats	airport	0	0	1	1
nordöstra	nordeastern	0	0	1	0
nordöstra	northeast	0	0	1	0
kritiskt	critical	0	0	1	0
ansökte	applied	0	0	1	0
instruktioner	instructions	0	0	1	1
mills	mills	0	0	1	0
fältet	the field	0	0	1	0
fältet	field	0	0	1	0
lindh	lindh	0	0	1	0
sinatra	sinatra	0	0	1	0
sekvens	sequence	0	0	1	1
kritiska	critical	0	0	1	0
best	best	0	0	1	0
linda	winding	0	0	1	0
linda	linda	0	0	1	0
viss	certain	0	0	1	1
viss	some	0	0	1	1
finsk	finnish	0	0	1	1
slutsatsen	concluded	0	0	1	0
slutsatsen	the conclusion	0	0	1	0
gävle	gävle	0	0	1	0
minoritet	minority	0	0	1	1
slovakien	slovakia	0	0	1	0
vardagen	the weekday	0	0	1	0
vardagen	everyday life	0	0	1	0
vardagen	vargaden	0	0	1	0
napoleons	napoleon's	0	0	1	0
napoleons	napoleon	0	0	1	0
visa	see	0	0	1	0
uppror	uprising	0	0	1	1
uppror	rebellion	0	0	1	1
guillou	guillou	0	0	1	0
medan	while	0	0	1	1
samhällets	society	0	0	1	0
samhällets	of society	0	0	1	0
synliga	visible	0	0	1	0
bred	broad	0	0	1	1
bokstaven	the letter	0	0	1	0
bokstaven	character	0	0	1	0
face	face	0	0	1	0
synligt	wisible	0	0	1	0
synligt	seen	0	0	1	0
synligt	visible	0	0	1	0
båt	boat	0	0	1	1
brev	letter	0	0	1	1
allmänheten	public	0	0	1	0
allmänheten	general public	0	0	1	0
beteende	behaviour	0	0	1	1
beteende	behavior	0	0	1	1
kärlek	love	0	0	1	1
mellanfot	metatarsus	1	1	0	0
mellanfot	metatarsal bones	1	1	0	0
mellanfot	metatarsel	1	0	1	0
mellanfot	metatarsals	1	0	1	0
mellanfot	metatarsal	1	1	0	0
mellanfot	mellanfot	1	0	1	0
mellanfot	islands	1	0	1	0
manchester	manchester	0	0	1	1
växande	growing	0	0	1	1
utmärkelser	commendations	0	0	1	0
utmärkelser	awards	0	0	1	0
rubrik	title	1	0	1	1
rubrik	headline	1	1	0	1
rubrik	many	1	0	1	0
rubrik	header	1	0	1	1
rubrik	quite a few	1	0	1	0
rubrik	riburk	1	0	1	0
rubrik	rubric	1	1	0	0
rubrik	runrik	1	0	1	0
rubrik	head line; rubric	1	0	1	0
rubrik	heading	1	0	1	1
bättre	better	0	0	1	1
hopp	hopes	0	0	1	0
hopp	hope	0	0	1	1
fursten	prince	0	0	1	0
sällskapshundar	pet dogs	0	0	1	0
sällskapshundar	companion dog	0	0	1	0
samisk	samian	0	0	1	0
samisk	sami	0	0	1	0
samisk	lapp	0	0	1	1
jan	jan	0	0	1	0
jan	january	0	0	1	0
utmärkelsen	award	0	0	1	0
utmärkelsen	the award	0	0	1	0
religionens	religion	0	0	1	0
religionens	religion's	0	0	1	0
liksom	and	0	0	1	0
liksom	as is	0	0	1	0
jah	jah	0	0	1	0
jag	i	0	0	1	1
ilska	anger	0	0	1	1
handla	act; buy; consume	0	0	1	0
handla	act	0	0	1	1
låna	borrow	0	0	1	1
låna	lana	0	0	1	0
lång	lang	0	0	1	0
lång	long	0	0	1	1
abba	abba	0	0	1	0
sociala	social	0	0	1	0
parlamentet	the parlament	0	0	1	0
parlamentet	parliament	0	0	1	0
fotbollsspelare	football player	0	0	1	0
fotbollsspelare	footballers	0	0	1	0
lucky	lucky	0	0	1	0
generalen	the general	0	0	1	0
generalen	general	0	0	1	0
bonde	bonde	0	0	1	0
bonde	farmer	0	0	1	1
parlamenten	parliaments	0	0	1	0
parlamenten	the parliament	0	0	1	0
traditionerna	traditions	0	0	1	0
traditionerna	the traditions	0	0	1	0
språk	language	0	0	1	1
meter	metre	0	0	1	1
meter	meters	0	0	1	0
meter	meter	0	0	1	1
underart	subspecies	0	0	1	0
tidigaste	earliest	0	0	1	0
tidigaste	tidigaste	0	0	1	0
britterna	british	0	0	1	0
britterna	the brits	0	0	1	0
omvärlden	world	0	0	1	0
omvärlden	surrounding world	0	0	1	0
omvärlden	outside world	0	0	1	0
h	h	0	0	1	0
rowling	rowling	0	0	1	0
effekterna	the effects	0	0	1	0
effekterna	effects	0	0	1	0
iranska	iranian	0	0	1	0
rymmer	has	0	0	1	0
rymmer	holds	0	0	1	0
premiärministern	the prime minister	0	0	1	0
premiärministern	prime minister	0	0	1	0
debuterade	debut	0	0	1	0
debuterade	debuted	0	0	1	0
koenigsegg	koenigsegg	0	0	1	0
michail	michail	0	0	1	0
priser	rates	0	0	1	0
priser	prizes	0	0	1	0
avlidit	perished	0	0	1	0
avlidit	died	0	0	1	0
priset	the prize	0	0	1	0
priset	rate	0	0	1	0
kronisk	chronic	0	0	1	1
minns	remembers	0	0	1	0
minns	remember	0	0	1	0
vietnams	vietnam	0	0	1	0
vietnams	vietnam's	0	0	1	0
mörkare	darkey	0	0	1	0
mörkare	darker	0	0	1	0
läkaren	the doctor	0	0	1	0
läkaren	physician	0	0	1	0
tvingade	forced	0	0	1	0
tvingade	forcing	0	0	1	0
populärkulturen	popular culture	0	0	1	0
förhållandena	conditions	0	0	1	0
förhållandena	the conditions	0	0	1	0
balansen	balance	0	0	1	0
balansen	the balance	0	0	1	0
kategorisvenskar	category swedes	0	0	1	0
undergång	during navigation	0	0	1	0
undergång	doom	0	0	1	1
undergång	destruction	0	0	1	1
striden	battle	0	0	1	0
striden	fight	0	0	1	0
finalen	final	0	0	1	0
bolivias	bolivia	0	0	1	0
bolivias	bolivia's	0	0	1	0
enda	only	0	0	1	1
enda	single	0	0	1	1
bilar	car	0	0	1	0
bilar	cars	0	0	1	0
ende	only	0	0	1	0
kedjor	chains	0	0	1	0
ett	a	0	0	1	1
ett	one; a; an	0	0	1	0
års	years	0	0	1	0
års	years (age)	0	0	1	0
års	year	0	0	1	0
marknaden	the market	0	0	1	0
marknaden	market	0	0	1	0
figuren	the character	0	0	1	0
figuren	figure	0	0	1	0
tycker	do	0	0	1	0
tycker	think	0	0	1	0
tycker	thinks	0	0	1	0
egypten	egypt	0	0	1	1
norge	norway	0	0	1	1
etc	etc.	0	0	1	0
harvard	harvard	0	0	1	0
marknader	markets	0	0	1	0
ogillade	disliked	0	0	1	0
ekvatorn	equator	0	0	1	0
ekvatorn	the equator	0	0	1	0
arbetat	worked	0	0	1	0
hårdrock	hard rock	0	0	1	0
hårdrock	hardrock	0	0	1	0
botten	the base	0	0	1	0
botten	bottom	0	0	1	1
co	co	0	0	1	0
co	coli	0	0	1	0
cm	centimeters	0	0	1	0
cm	cm	0	0	1	0
cc	cc	0	0	1	0
malcolm	malcolm	0	0	1	0
mengele	mengele	0	0	1	0
cd	cd	0	0	1	0
sannolikhet	probability	0	0	1	1
stabila	stable	0	0	1	0
musikvideo	music video	0	0	1	0
cp	cp	0	0	1	0
gudarnas	the gods'	0	0	1	0
gudarnas	gods	0	0	1	0
gudarnas	god's	0	0	1	0
utlöste	triggered	0	0	1	0
antal	number of	0	0	1	0
antal	number	0	0	1	1
jussi	jussi	0	0	1	0
keltiska	celtic	0	0	1	1
moraliskt	morally	0	0	1	1
moraliskt	moralist	0	0	1	0
moraliskt	moral	0	0	1	0
högskolor	colleges	0	0	1	0
högskolor	hogskoñor	0	0	1	0
centralort	central city	0	0	1	0
centralort	regional centre	0	0	1	0
centralort	centralot	0	0	1	0
rockband	rock band	0	0	1	0
genetik	genetics	0	0	1	1
förlusterna	the losses	0	0	1	0
förlusterna	loss	0	0	1	0
louisiana	louisiana	0	0	1	0
antas	is required	0	0	1	0
antas	assumed	0	0	1	0
antas	expected (to)	0	0	1	0
antar	adopting	0	0	1	0
antar	adopt	0	0	1	0
antar	suppose	0	0	1	0
typisk	typical	0	0	1	1
molekyler	molecules	0	0	1	0
lägenhet	apartment	0	0	1	1
lägenhet	appartment	0	0	1	0
upplösningen	dissolution	0	0	1	0
upplösningen	disbandment	0	0	1	0
lämpligt	suitable	0	0	1	0
lämpligt	fitness	0	0	1	0
berättelse	tale	0	0	1	1
berättelse	story	0	0	1	1
berättelse	's re	0	0	1	0
lämpliga	suitable	0	0	1	0
råolja	crude oil	0	0	1	1
hänvisade	referenced	0	0	1	0
hänvisade	refer	0	0	1	0
hänvisade	referred	0	0	1	0
lägger	put	0	0	1	0
lägger	lies	0	0	1	0
lägger	add	0	0	1	0
mandatperiod	term	0	0	1	0
mandatperiod	term (of office)	0	0	1	0
mandatperiod	term of office	0	0	1	0
tjorven	tjorven	0	0	1	0
weber	weber	0	0	1	0
rikets	its	0	0	1	0
rikets	the kingdom's	0	0	1	0
rikets	the realms	0	0	1	0
demokrati	democracy	0	0	1	1
aktivitet	activity	0	0	1	1
installera	installing	0	0	1	0
installera	install	0	0	1	1
vd	ceo	0	0	1	0
ondskan	the evil	0	0	1	0
ondskan	evil	0	0	1	0
vi	we	0	0	1	1
ryssland	russia	0	0	1	1
site	site	0	0	1	0
längst	farthest	0	0	1	1
längst	longest	0	0	1	0
längst	at	0	0	1	0
lust	desire	0	0	1	1
lust	loss	0	0	1	0
vs	vs	0	0	1	0
flickor	girls	0	0	1	0
skapare	creator	0	0	1	1
säkerhetspolitik	safety policy	0	0	1	0
säkerhetspolitik	security	0	0	1	0
säkerhetspolitik	security policy	0	0	1	0
sitt	his	0	0	1	1
sitt	its	0	0	1	0
slovenska	slovenian	0	0	1	0
sysselsätter	employs	0	0	1	0
evenemang	event	0	0	1	1
nobelkommittén	the nobel commitee	0	0	1	0
tupac	tupac	0	0	1	0
juan	juan	0	0	1	0
juan	mr juan	0	0	1	0
medeltida	middleaged	0	0	1	0
medeltida	medival	0	0	1	0
medeltida	medieval	0	0	1	1
foundationthe	foundationthe	0	0	1	0
foundationthe	the foundation	0	0	1	0
huden	skin	0	0	1	0
romance	romance	0	0	1	0
matthew	matthew	0	0	1	0
färg	colors	0	0	1	0
färg	colour	0	0	1	1
terrorism	terrorism	0	0	1	1
flesta	most	0	0	1	1
ball	ball	0	0	1	0
columbia	columbia	0	0	1	0
columbia	colombia	0	0	1	0
sade	said	0	0	1	0
tävlingar	competitions	0	0	1	0
tävlingar	contests	0	0	1	0
konstantin	konstantin	0	0	1	0
konstantin	constantine	0	0	1	0
nederlag	defeat	0	0	1	1
anfield	anfield	0	0	1	0
ikea	ikea	0	0	1	0
sjukhus	hospital	0	0	1	1
sjukhus	hospitals	0	0	1	0
knäppupp	knäppup	0	0	1	0
knäppupp	knäppupp	0	0	1	0
diabetes	diabetes	0	0	1	1
isländska	icelandic	0	0	1	0
lupus	lupus	0	0	1	1
off	off	0	0	1	0
ledde	resulted	0	0	1	0
ledde	led	0	0	1	0
ledda	led	0	0	1	0
ledda	run (by)	0	0	1	0
versaillesfreden	versailles peace	0	0	1	0
versaillesfreden	treaty of versailles	0	0	1	0
lägre	lower	0	0	1	1
gatan	street	0	0	1	0
gatan	the street	0	0	1	0
kontakt	plug	0	0	1	0
kontakt	contact	0	0	1	1
paus	pause	0	0	1	1
paus	paus	0	0	1	0
aktuell	current	0	0	1	1
kvast	broom	1	1	0	1
kvast	factories	1	0	1	0
kvast	groom	1	0	1	0
köpenhamns	kopenhamns	0	0	1	0
köpenhamns	copenhagen	0	0	1	0
köpenhamns	copenhagen's	0	0	1	0
ståndpunkt	standpoint	0	0	1	1
ståndpunkt	position	0	0	1	0
paul	paul	0	0	1	0
flest	most	0	0	1	0
flest	the most	0	0	1	0
tolkade	interpreted	0	0	1	0
derivata	derivative	0	0	1	0
kunder	customer	0	0	1	0
kunder	customers	0	0	1	0
kunder	clients	0	0	1	0
nacional	nacional	0	0	1	0
englands	england's	0	0	1	0
planeten	planet	0	0	1	0
planeten	the planet	0	0	1	0
kosovos	kosovo	0	0	1	0
kosovos	kosovo's	0	0	1	0
filmens	the film's	0	0	1	0
filmens	film	0	0	1	0
framtid	future	0	0	1	1
gärningar	yarn penetrations	0	0	1	0
gärningar	deeds	0	0	1	0
government	government	0	0	1	0
ledarna	the leaders	0	0	1	0
ledarna	conductors	0	0	1	0
grönwall	gronwall	0	0	1	0
grönwall	grönwall	0	0	1	0
arbetarklassen	working class	0	0	1	0
arbetarklassen	the working class	0	0	1	0
halvön	peninsula	0	0	1	0
halvön	the peninsula	0	0	1	0
pressas	pressed	0	0	1	0
karaktär	character	0	0	1	1
insåg	realized	0	0	1	0
emma	emaa	0	0	1	0
emma	emma	0	0	1	0
aktiebolag	companies	0	0	1	0
aktiebolag	stock company	0	0	1	0
aktiebolag	limited company; joint-stock company	0	0	1	0
vallhund	herder	0	0	1	0
vallhund	herding dog	0	0	1	0
stadsbild	cityscape	0	0	1	1
amazonas	the amazon rainforest	0	0	1	0
amazonas	amazon	0	0	1	0
amazonas	amazonas	0	0	1	0
symptomen	symptoms	0	0	1	0
symptomen	the symptoms	0	0	1	0
därtill	thereto	0	0	1	1
flotta	fleet	0	0	1	1
järnmalm	iron ore	0	0	1	0
järnmalm	jarnmalm	0	0	1	0
tackade	thanked	0	0	1	0
tackade	said/thanked	0	0	1	0
bredare	wider	0	0	1	1
bredare	broad	0	0	1	0
miniatyr|	miniature	0	0	1	0
filmografi	filmography	0	0	1	0
filmografi	folmografi	0	0	1	0
anarkismen	the anarkism	0	0	1	0
anarkismen	anarchism	0	0	1	0
trotskij	trotskij	0	0	1	0
trotskij	trotsky	0	0	1	0
vägar	roads	0	0	1	0
vägar	paths	0	0	1	0
avstånd	distance	0	0	1	1
stannar	stay	0	0	1	0
stannar	stop	0	0	1	0
stannar	stays	0	0	1	0
föreställningar	performances	0	0	1	0
föreställningar	notions	0	0	1	0
transport	carriage	0	0	1	1
transport	transportation	0	0	1	1
transport	transport	0	0	1	1
skriftliga	written	0	0	1	0
atomkärnor	nuclei	0	0	1	0
atomkärnor	nuclear particles	0	0	1	0
atomkärnor	atomic cores	0	0	1	0
påvisa	detection	0	0	1	0
påvisa	prove	0	0	1	1
påvisa	show	0	0	1	1
februari	february	0	0	1	1
februari	februari	0	0	1	0
kolonin	colony	0	0	1	0
behandlades	treated	0	0	1	0
flitigt	actively	0	0	1	0
flitigt	frequent	0	0	1	0
dags	time	0	0	1	0
försäkra	insure	0	0	1	1
försäkra	make sure	0	0	1	0
försäkra	assure	0	0	1	1
naturlig	natural	0	0	1	1
kollektivtrafik	public transport	0	0	1	0
begränsas	limited	0	0	1	0
begränsas	(gets) limited	0	0	1	0
begränsas	begransas	0	0	1	0
begränsar	limit	0	0	1	0
begränsar	limits	0	0	1	0
ateist	atheist	0	0	1	1
svaga	faint	0	0	1	0
svaga	weak	0	0	1	0
begränsat	limited	0	0	1	0
begränsat	restricted	0	0	1	0
mönster	marks	0	0	1	0
halland	halland	0	0	1	0
svagt	weak	0	0	1	0
gandalf	gandalf	0	0	1	0
vargen	the wolf	0	0	1	0
lär	teach	0	0	1	0
lär	learn	0	0	1	0
begränsad	restricted	0	0	1	0
begränsad	limited	0	0	1	1
jämföras	comparable	0	0	1	0
jämföras	compared	0	0	1	0
kontinenten	the continent	0	0	1	0
blodiga	blooded	0	0	1	0
blodiga	bloody	0	0	1	0
angeles	angeles	0	0	1	0
försvann	disappeared	0	0	1	0
kontinenter	continents	0	0	1	0
warner	warner	0	0	1	0
absint	absinthe	0	0	1	0
hittills	date	0	0	1	0
hittills	so far	0	0	1	0
burma	burma	0	0	1	1
anpassade	adjusted	0	0	1	0
anpassade	custom	0	0	1	0
sekelskiftet	turn	0	0	1	0
sekelskiftet	the turn of the century	0	0	1	0
planetens	planet	0	0	1	0
planetens	the planets	0	0	1	0
kristus	christ	0	0	1	1
lund	grove	0	0	1	1
lund	lund	0	0	1	0
mera	more	0	0	1	1
gräslök	chive	1	0	1	1
gräslök	culture	1	0	1	0
gräslök	chives	1	1	0	0
gräslök	raslok	1	0	1	0
varma	hot	0	0	1	0
varma	warm	0	0	1	0
päls	fur	0	0	1	1
nåd	mercy	0	0	1	0
nåd	grace	0	0	1	1
peters	peters	0	0	1	0
skola	school	0	0	1	1
missnöjet	discontent	0	0	1	0
missnöjet	grievance	0	0	1	0
hudfärg	color	0	0	1	0
hudfärg	skin color	0	0	1	0
når	reach	0	0	1	0
når	when	0	0	1	0
når	reaches	0	0	1	0
nås	nas	0	0	1	0
nås	is reached	0	0	1	0
nås	reached	0	0	1	0
tina	defrost	0	0	1	0
tina	thaw	0	0	1	1
tina	tina	0	0	1	0
radioaktiva	radioactive	0	0	1	0
samlingar	collections	0	0	1	0
samlingar	collection	0	0	1	0
uppvisade	showed	0	0	1	0
indonesien	indonesia	0	0	1	1
apollo	apollo	0	0	1	0
radioaktivt	radioactive	0	0	1	0
öppnades	were opened	0	0	1	0
öppnades	was opened	0	0	1	0
öppnades	opened	0	0	1	0
lättare	light	0	0	1	0
lättare	easier	0	0	1	0
official	official	0	0	1	0
volvo	volvo	0	0	1	0
ruset	ruset	0	0	1	0
ruset	the fuddle	0	0	1	0
ruset	intoxication	0	0	1	0
stormakt	great power	0	0	1	1
stormakt	major power	0	0	1	0
monument	monuments	0	0	1	0
monument	monument	0	0	1	1
distribution	distribution	0	0	1	1
baptism	baptist	1	1	0	0
baptism	bapist faith	1	1	0	0
baptism	baptist faith	1	1	0	1
baptism	universe	1	0	1	0
baptism	döpare	1	0	1	0
baptism	the universe	1	0	1	0
baptism	baptists	1	1	0	0
baptism	baptism	1	1	0	0
butiker	shops	0	0	1	0
butiker	stores	0	0	1	0
närmar	close	0	0	1	0
närmar	closing	0	0	1	0
närmar	close in	0	0	1	0
möjliggör	enable	0	0	1	0
möjliggör	enables	0	0	1	0
leukemi	leukemia	0	0	1	1
självklart	course	0	0	1	0
heter	units	0	0	1	0
heter	is named	0	0	1	0
heter	(is the) name (of)	0	0	1	0
utnyttjar	using	0	0	1	0
utnyttjar	uses	0	0	1	0
utnyttjas	utilized	0	0	1	0
utnyttjas	used	0	0	1	0
separerade	separated	0	0	1	0
fågel	bird	0	0	1	1
broder	brother	0	0	1	1
banan	the track	0	0	1	0
banan	banana	0	0	1	1
vitryssland	belarus	0	0	1	0
sharia	sharia	0	0	1	0
programmet	program	0	0	1	0
programmet	the application	0	0	1	0
programmet	the program	0	0	1	0
brandenburg	brandenburg	0	0	1	0
distinkta	distinct	0	0	1	0
lutning	closing	0	0	1	0
lutning	angle	0	0	1	0
lutning	incline	0	0	1	1
relationen	the relation	0	0	1	0
relationen	ratio	0	0	1	0
oavgjort	tie	0	0	1	0
oavgjort	draw	0	0	1	0
modernistiska	modernistic	0	0	1	0
modernistiska	modernist	0	0	1	0
köpte	purchased	0	0	1	0
köpte	bought	0	0	1	0
francisco	francisco	0	0	1	0
francisco	fransisco	0	0	1	0
uttalade	commented; made a comment; spoke about	0	0	1	0
uttalade	spoke	0	0	1	0
uttalade	stated	0	0	1	0
tider	times; ages	0	0	1	0
tider	times	0	0	1	0
söner	sons	0	0	1	0
tiden	the time	0	0	1	0
tiden	time	0	0	1	0
hård	diffcult	0	0	1	0
hård	hard	0	0	1	1
inspiration	inspiration	0	0	1	1
syskon	sibling	0	0	1	1
syskon	siblings	0	0	1	0
mozart	mozart	0	0	1	0
mineraler	minerals	0	0	1	0
provinser	provinces	0	0	1	0
resulterade	resulted	0	0	1	0
rötter	roots	0	0	1	0
brevet	the letter	0	0	1	0
brevet	letter	0	0	1	0
child	child	0	0	1	0
elisabeth	elisabeth	0	0	1	0
glädje	joy	0	0	1	1
områdets	the area's	0	0	1	0
områdets	of the area	0	0	1	0
områdets	area	0	0	1	0
bosniska	bosnian	0	0	1	0
representanthuset	house of representatives	0	0	1	1
invadera	invade	0	0	1	1
preussen	prussia	0	0	1	1
konsekvenserna	impact	0	0	1	0
konsekvenserna	consequensis	0	0	1	0
barmel	barmel	0	0	1	0
bibel	bible	0	0	1	1
bibel	insulin	0	0	1	0
bibel	bilble	0	0	1	0
spel	game	0	0	1	1
edward	edward	0	0	1	0
grundande	founding	0	0	1	0
spannmål	cereals	0	0	1	1
spannmål	grain	0	0	1	1
brushane	secondary	1	0	1	0
brushane	rushane	1	0	1	0
brushane	bird	1	1	0	0
brushane	brushane (bird)	1	0	1	0
brushane	ruff	1	1	0	1
ale	ale	0	0	1	0
längd	length	0	0	1	1
parterna	parties	0	0	1	0
golvet	the floor	0	0	1	0
golvet	floor	0	0	1	0
tjäna	profit	0	0	1	0
tjäna	earn	0	0	1	1
tjäna	make	0	0	1	1
längs	along	0	0	1	1
vidsträckta	broad	0	0	1	0
vidsträckta	wide; broad	0	0	1	0
geologi	geology	0	0	1	1
jacob	jacob	0	0	1	0
skolor	schools	0	0	1	0
föder	give birth	0	0	1	0
föder	give birth of	0	0	1	0
föder	gives birth	0	0	1	0
innefattar	comprises	0	0	1	0
innefattar	includes	0	0	1	0
uttryck	expression	0	0	1	1
målning	painting	0	0	1	1
bipolär	bipolar	0	0	1	1
upplöstes	dissolved	0	0	1	0
estland	estland	0	0	1	0
estland	estonia	0	0	1	1
jamaica	jamaica	0	0	1	1
starkast	strongest	0	0	1	0
vänstern	the left wing	0	0	1	0
vänstern	left party	0	0	1	0
vänstern	western	0	0	1	0
galax	galaxy	0	0	1	1
horn	horn	0	0	1	1
horn	horns	0	0	1	0
chef	head	0	0	1	1
alltsedan	even since	0	0	1	0
alltsedan	since	0	0	1	1
eurovision	eurovision	0	0	1	0
renässans	renaissance	0	0	1	1
italiens	italy's	0	0	1	0
italiens	italian	0	0	1	0
verksamma	active	0	0	1	0
kraftfull	forceful	0	0	1	1
kraftfull	powerful	0	0	1	1
speglar	mirrors	0	0	1	0
speglar	mirror	0	0	1	0
tolv	twelve	0	0	1	1
stadskärna	town	0	0	1	0
stadskärna	city core	0	0	1	0
stadskärna	town centre	0	0	1	0
stadskärna	city center	0	0	1	0
vampyr	vampire	0	0	1	1
cyklar	bicycles	0	0	1	0
cyklar	bikes	0	0	1	0
cyklar	cycles	0	0	1	0
mellanöstern	middle	0	0	1	0
mellanöstern	the middle east	0	0	1	0
mellanöstern	middle east	0	0	1	0
hovrätten	court of appeals	0	0	1	0
hovrätten	the court of appeal	0	0	1	0
bidrar	contributes	0	0	1	0
petra	petra	0	0	1	0
musikalen	the musical	0	0	1	0
griffin	griffin	0	0	1	0
innanför	inside	0	0	1	1
innanför	within	0	0	1	1
pluto	pluto	0	0	1	1
rapporterar	reports	0	0	1	0
norstedt	norstedt	0	0	1	0
olsson	olsson	0	0	1	0
studeras	studied	0	0	1	0
studeras	(is) studied	0	0	1	0
studeras	is studied	0	0	1	0
sidan	page	0	0	1	0
sidan	the side	0	0	1	0
sidan	side	0	0	1	0
regerande	reigning	0	0	1	0
regerande	ruling	0	0	1	1
stoft	dust	0	0	1	1
månader	months	0	0	1	0
placerades	placed	0	0	1	0
månaden	the month	0	0	1	0
månaden	months	0	0	1	0
månaden	month	0	0	1	0
akc	akc	0	0	1	0
lön	salary	0	0	1	1
lön	wage; salary	0	0	1	0
melankoli	melancholy	0	0	1	1
kongressen	congress	0	0	1	0
faktiskt	in fact; actually; indeed	0	0	1	0
faktiskt	actually	0	0	1	1
faktiskt	really	0	0	1	1
bro	bridge	0	0	1	1
tillsammans	together	0	0	1	1
föreställer	picture	0	0	1	0
föreställer	depicts	0	0	1	0
föreställer	pictures	0	0	1	0
faktiska	actual	0	0	1	0
total	total	0	0	1	1
absolution	absolution	0	0	1	1
sarah	sarah	0	0	1	0
ställas	set	0	0	1	0
ställas	be set	0	0	1	0
ställas	prepared	0	0	1	0
negativa	negative	0	0	1	0
karaktärer	character	0	0	1	0
karaktärer	characters	0	0	1	0
karaktären	the character	0	0	1	0
karaktären	character	0	0	1	0
utfördes	carried out	0	0	1	0
utfördes	was carried out	0	0	1	0
utfördes	preformed	0	0	1	0
indiana	indiana	0	0	1	0
tempererat	temperate	0	0	1	0
tempererat	tempered	0	0	1	0
negativt	negative	0	0	1	0
supportrar	supports	0	0	1	0
supportrar	supporters	0	0	1	0
ifall	if	0	0	1	1
genomför	implement	0	0	1	0
genomför	carry out	0	0	1	0
genomför	out	0	0	1	0
giovanni	giovanni	0	0	1	0
fingrar	finger	0	0	1	0
fingrar	fingers	0	0	1	0
award	award	0	0	1	0
sydöstra	the southeast	0	0	1	0
sydöstra	south east	0	0	1	0
sydöstra	south eastern	0	0	1	0
åtminstone	at least	0	0	1	1
nku	nku	0	0	1	0
synsätt	effects	0	0	1	0
synsätt	viewpoint	0	0	1	0
synsätt	effect	0	0	1	0
alces	alces	0	0	1	0
bemärkelse	meaning	0	0	1	0
bemärkelse	sense	0	0	1	1
springer	running	0	0	1	0
springer	springer	0	0	1	0
absorberas	absorbed	0	0	1	0
absorberas	(gets) absorbed	0	0	1	0
friheten	freedom; liberty	0	0	1	0
friheten	freedom	0	0	1	0
friheten	liberty	0	0	1	0
ik	ik	0	0	1	0
förlängning	overtime; extension; prolongation	0	0	1	0
förlängning	extension	0	0	1	1
era	era	0	0	1	1
era	yours	0	0	1	0
transparency	transparency	0	0	1	0
zirkon	assisted	1	0	1	0
zirkon	contributed	1	0	1	0
zirkon	zirconium	1	1	0	0
zirkon	zircon	1	1	0	0
zirkon	zirkon	1	1	0	0
zirkon	further	1	0	1	0
föregångaren	predecessor	0	0	1	0
föregångaren	it's predecessor	0	0	1	0
skiljer	differs	0	0	1	0
skiljer	is different; differ	0	0	1	0
skiljer	different	0	0	1	0
vietnamesiska	vietnamese	0	0	1	0
gloria	gloria	0	0	1	0
vackra	beautiful	0	0	1	0
vackra	fine	0	0	1	0
felaktiga	false	0	0	1	0
ekonomiskt	economic	0	0	1	0
ekonomiskt	economically	0	0	1	1
ekonomiskt	economical	0	0	1	0
sommar	summer	0	0	1	1
indien	india	0	0	1	1
felaktigt	incorrect	0	0	1	0
felaktigt	erronenous	0	0	1	0
felaktigt	error	0	0	1	0
indier	indians	0	0	1	0
enhet	unit	0	0	1	1
enhet	entity	0	0	1	1
valborg	may day	0	0	1	0
valborg	valborg	0	0	1	0
förenta	united	0	0	1	0
utlandet	foreign land	0	0	1	0
utlandet	abroad	0	0	1	0
utlandet	foreign	0	0	1	0
gotlands	gotland's	0	0	1	0
gotlands	gotland	0	0	1	0
ansluter	connects	0	0	1	0
ansluter	connect	0	0	1	0
protestantiska	protestant	0	0	1	0
protestantiska	protestantic	0	0	1	0
firar	celebrates	0	0	1	0
firar	celebrate	0	0	1	0
gillar	like	0	0	1	0
gillar	enjoy; like	0	0	1	0
gillar	likes	0	0	1	0
övergrepp	assault	0	0	1	0
övergrepp	abuse	0	0	1	0
övergrepp	assult (-s)	0	0	1	0
beach	beach	0	0	1	0
sammansatt	composed	0	0	1	0
sammansatt	compound	0	0	1	1
mötet	the meeting	0	0	1	0
mötet	meeting	0	0	1	0
biografer	movie theaters	0	0	1	0
biografer	movie theaters; cinemas	0	0	1	0
biografer	cinemas	0	0	1	0
möter	meet	0	0	1	0
möter	meets	0	0	1	0
kategorieuropas	category europe	0	0	1	0
lag	law	0	0	1	1
lag	act	0	0	1	1
koreakriget	korean war	0	0	1	0
koreakriget	the korean war	0	0	1	0
davis	davis	0	0	1	0
visste	did	0	0	1	0
lat	methacrylate	0	0	1	0
höjdpunkt	highlight	0	0	1	0
höjdpunkt	climax	0	0	1	1
höjdpunkt	high point	0	0	1	0
möten	moten	0	0	1	0
möten	meetings	0	0	1	0
orden	the words	0	0	1	0
orden	words	0	0	1	0
medlemsstat	member state	0	0	1	0
green	green	0	0	1	0
massmedia	media	0	0	1	0
massmedia	mass media	0	0	1	1
livets	life's	0	0	1	0
livets	life	0	0	1	0
livets	the life's	0	0	1	0
ordet	the word	0	0	1	0
ordet	word	0	0	1	0
order	order	0	0	1	1
order	words	0	0	1	0
förhistoria	prehistory	0	0	1	1
natten	overnight	0	0	1	0
office	office	0	0	1	0
förkortning	abbreviation	0	0	1	1
alltför	all too	0	0	1	0
alltför	exessive	0	0	1	0
alltför	way too	0	0	1	0
exempel	example	0	0	1	1
exempel	for example; for instance; sample(-s)	0	0	1	0
ramadan	ramadan	0	0	1	0
blandning	mix	0	0	1	1
blandning	mixture	0	0	1	1
japan	japan	0	0	1	1
bidra	contribute	0	0	1	0
världen	world	0	0	1	0
världen	the world	0	0	1	0
lösas	solved	0	0	1	0
straff	penalty	0	0	1	1
straff	punishment	0	0	1	1
straff	punishments	0	0	1	0
lagets	the team's	0	0	1	0
lagets	substrate	0	0	1	0
frågor	questions	0	0	1	0
väljs	selected	0	0	1	0
väljs	elect	0	0	1	0
fragment	fragment	0	0	1	1
fragment	fragments	0	0	1	0
vanligtvis	usually	0	0	1	1
vanligtvis	generally	0	0	1	0
främsta	primary; foremost; primarily; principally	0	0	1	0
främsta	request	0	0	1	0
främsta	primary	0	0	1	0
främste	chief	0	0	1	0
främste	premier	0	0	1	0
kategoriledamöter	category members	0	0	1	0
kategoriledamöter	category: members	0	0	1	0
band	band	0	0	1	1
band	tape	0	0	1	1
fredsbevarande	fresberarande	0	0	1	0
fredsbevarande	peace	0	0	1	0
fredsbevarande	peacekeeping	0	0	1	0
bana	course	0	0	1	1
bana	web	0	0	1	0
they	they	0	0	1	0
spelningen	the gig	0	0	1	0
spelningen	the concert	0	0	1	0
rättsliga	justice	0	0	1	0
rättsliga	legal	0	0	1	0
bank	bank	0	0	1	1
genomförts	out	0	0	1	0
stående	standing	0	0	1	1
stående	above	0	0	1	0
ansvariga	charge	0	0	1	0
huvudartikel	main article	0	0	1	0
huvudartikel	principal article	0	0	1	0
helvetet	hell	0	0	1	0
helvetet	the hell	0	0	1	0
l	l	0	0	1	0
grannar	neighbors	0	0	1	1
grannar	neighbours	0	0	1	1
diskuteras	discussed	0	0	1	0
diskuteras	is discucssed	0	0	1	0
knutpunkt	hub	0	0	1	0
tendens	tendency	0	0	1	1
föreslogs	suggested	0	0	1	0
föreslogs	was suggested	0	0	1	0
föreslogs	proposed	0	0	1	0
carlos	carlos	0	0	1	0
tillgängligt	available	0	0	1	0
germanska	germanic	0	0	1	0
germanska	germanian	0	0	1	0
inflytandet	the influence	0	0	1	0
inflytandet	inflytandet	0	0	1	0
inflytandet	influence	0	0	1	0
moçambique	mozambique	0	0	1	0
koldioxid	carbon dioxide	0	0	1	1
koldioxid	co	0	0	1	0
tillgängliga	available	0	0	1	0
voddler	voddler	0	0	1	0
framställa	represent; depict; produce	0	0	1	0
framställa	produce	0	0	1	1
framställa	the installation	0	0	1	0
trädde	met	0	0	1	0
trädde	entered	0	0	1	0
trädde	come into effect	0	0	1	0
kejserliga	imperially	0	0	1	0
kejserliga	imperial	0	0	1	0
framställs	is depicted	0	0	1	0
framställs	prepared	0	0	1	0
daniel	daniel	0	0	1	0
trafik	traffic	0	0	1	1
bruttonationalprodukt	gross national product	0	0	1	0
bruttonationalprodukt	gross domestic product	0	0	1	0
bruttonationalprodukt	bnp	0	0	1	0
oskar	oskar	0	0	1	0
vete	wheat	0	0	1	1
klimatet	environment	0	0	1	0
klimatet	climate	0	0	1	0
klimatet	the climate	0	0	1	0
öknen	the desert	0	0	1	0
öknen	desert	0	0	1	0
veta	know	0	0	1	1
veta	out	0	0	1	0
sedermera	subsequently	0	0	1	0
sedermera	since	0	0	1	1
veto	veto	0	0	1	1
veto	vetoe	0	0	1	0
standard	standard	0	0	1	1
tillbaka	back	0	0	1	1
upprättandet	establishment	0	0	1	0
upprättandet	establishing	0	0	1	0
förmögenhet	fortune	0	0	1	1
förmögenhet	wealth	0	0	1	0
vågade	dared	0	0	1	0
ange	set	0	0	1	0
ange	name	0	0	1	0
sprit	liqeur	0	0	1	0
sprit	alcohol	0	0	1	1
förblev	remained	0	0	1	1
professionell	professional	0	0	1	1
fåtal	few	0	0	1	0
fåtal	a few	0	0	1	0
sändas	broadcast	0	0	1	0
sändas	be transmitted	0	0	1	0
sändas	sent	0	0	1	0
personerna	people; persons	0	0	1	0
personerna	subjects	0	0	1	0
personerna	the persons	0	0	1	0
öst	east	0	0	1	1
hänvisar	reference	0	0	1	0
möjlig	possible	0	0	1	1
another	another	0	0	1	0
statskupp	coup	0	0	1	0
ingmar	ingmar	0	0	1	0
synnerligen	remarkably; particularly	0	0	1	0
synnerligen	particularly	0	0	1	1
synnerligen	quite	0	0	1	0
drabbade	suffering	0	0	1	0
drabbade	affected	0	0	1	0
är	is	0	0	1	0
ingen	there is no	0	0	1	0
ingen	no	0	0	1	1
lidande	sufferer	0	0	1	0
inget	not	0	0	1	0
inget	no	0	0	1	0
john	john	0	0	1	0
dogs	dogs	0	0	1	0
medborgare	citizens	0	0	1	0
antisemitismen	antisemitism	0	0	1	0
antisemitismen	anti-semitism	0	0	1	0
albert	albert	0	0	1	0
kvarvarande	remaining	0	0	1	1
kvarvarande	residual	0	0	1	0
kvarvarande	lasting	0	0	1	0
persson	persson	0	0	1	0
bojkott	boycott	0	0	1	1
kraftverk	plant	0	0	1	0
kraftverk	power plant	0	0	1	1
trupp	troop	0	0	1	1
trupp	troops	0	0	1	0
kände	felt	0	0	1	0
zeeland	zealand	0	0	1	0
zeeland	zeeland	0	0	1	0
omröstningen	vote	0	0	1	0
omröstningen	the election	0	0	1	0
religionerna	religions	0	0	1	0
religionerna	the religions	0	0	1	0
toronto	toronto	0	0	1	0
binda	bind	0	0	1	1
binda	tying	0	0	1	0
binda	bond	0	0	1	0
kronan	swedish krona	0	0	1	0
kronan	crown	0	0	1	0
kronan	kronan	0	0	1	0
sonen	the son	0	0	1	0
scener	scenes	0	0	1	0
scenen	the stage	0	0	1	0
scenen	stage	0	0	1	0
binds	bind	0	0	1	0
binds	bound	0	0	1	0
binds	(is) bound	0	0	1	0
tjänsten	the service	0	0	1	0
tjänsten	service	0	0	1	0
iron	iron	0	0	1	1
byggts	built	0	0	1	0
minut	minute	0	0	1	1
pelle	pellet	0	0	1	0
pelle	pelle	0	0	1	0
utsläpp	emission	0	0	1	0
utsläpp	emissions	0	0	1	0
värsta	worst	0	0	1	0
skolorna	schools	0	0	1	0
skolorna	the schools	0	0	1	0
mannen	art	0	0	1	0
mannen	the man	0	0	1	0
onani	masturbation	0	0	1	1
münchen	munchen	0	0	1	0
münchen	munich	0	0	1	0
åke	åke	0	0	1	0
göring	goring	0	0	1	0
göring	cleaning	0	0	1	0
omvandling	transformation	0	0	1	1
framtida	future	0	0	1	1
koloniala	colonial	0	0	1	0
anledningar	reasons	0	0	1	0
kalendern	calendar	0	0	1	0
kalendern	calender	0	0	1	0
stavning	spelling	0	0	1	1
magnus	magnus	0	0	1	0
aftonbladet	aftonbladet	0	0	1	0
aftonbladet	newsweek	0	0	1	0
aftonbladet	the evening paper	0	0	1	0
lades	put	0	0	1	0
lades	was	0	0	1	0
figurerna	figures	0	0	1	0
figurerna	characters	0	0	1	0
verkat	worked	0	0	1	0
verkat	acted	0	0	1	0
verkat	seemed	0	0	1	0
verkar	acting	0	0	1	0
verkar	seems	0	0	1	0
verkar	operates	0	0	1	0
maiden	maiden	0	0	1	0
bruce	bruce	0	0	1	0
värdet	the value	0	0	1	0
stödja	support	0	0	1	1
what	what	0	0	1	0
skansen	forecastle	0	0	1	0
värden	values	0	0	1	0
hälften	the one half	0	0	1	0
hälften	half	0	0	1	0
verkan	effect	0	0	1	1
flygplatsen	airport	0	0	1	0
flygplatsen	the airport	0	0	1	0
årens	the year's	0	0	1	0
årens	years	0	0	1	0
aminosyra	amino acid	0	0	1	1
eviga	eternal	0	0	1	0
freja	freja	0	0	1	0
freja	joe	0	0	1	0
bortom	beyond	0	0	1	1
bortom	beyond the	0	0	1	0
sammanhängande	connective	0	0	1	0
sammanhängande	context of	0	0	1	0
sammanhängande	continous	0	0	1	0
evigt	forever	0	0	1	1
evigt	eternal	0	0	1	0
åskådare	spectators	0	0	1	0
åskådare	audience; viewer	0	0	1	0
gräns	border	0	0	1	1
gräns	limit	0	0	1	1
effekten	the effect	0	0	1	0
effekten	effect	0	0	1	0
män	males	0	0	1	0
män	men	0	0	1	0
mitten	middle	0	0	1	1
mitten	mid	0	0	1	0
damer	ladies	0	0	1	0
glödlampor	lightbulbs	0	0	1	0
glödlampor	light bulbs	0	0	1	0
glödlampor	filament	0	0	1	0
lewis	lewis	0	0	1	0
turnén	turn	0	0	1	0
turnén	tour	0	0	1	0
turnén	tournament	0	0	1	0
hinduiska	hindu	0	0	1	0
biträdande	assistant	0	0	1	1
biträdande	assisting	0	0	1	0
biträdande	deputy	0	0	1	0
madeira	madeira	0	0	1	1
effekter	effeckter	0	0	1	0
effekter	effects; repercussions	0	0	1	0
effekter	effects	0	0	1	0
capitol	capitol	0	0	1	0
rankning	ranking	0	0	1	0
rankning	rating	0	0	1	0
någonstans	somewhere	0	0	1	1
någonstans	nowhere	0	0	1	0
estetiska	aesthetic	0	0	1	0
arthur	arthur	0	0	1	0
ambassad	embassy	0	0	1	1
välstånd	prosperity	0	0	1	1
välstånd	salstand	0	0	1	0
kejsar	emperor	0	0	1	0
variera	vary	0	0	1	1
försämrades	worsened	0	0	1	0
försämrades	worsening	0	0	1	0
försämrades	decreased	0	0	1	0
namn	name	0	0	1	1
kontinuerlig	continuous	0	0	1	1
imperium	empire	0	0	1	1
dj	dj	0	0	1	0
di	di	0	0	1	0
motstånd	resistance	0	0	1	1
motstånd	opposition	0	0	1	1
de	the	0	0	1	1
de	they	0	0	1	1
dc	d.c.	0	0	1	0
da	da	0	0	1	0
stalins	stalins	0	0	1	0
stalins	stalin	0	0	1	0
watson	watson	0	0	1	0
orolig	worried	0	0	1	1
riktningen	direction	0	0	1	0
riktningen	denomination	0	0	1	0
ändra	change	0	0	1	1
du	to	0	0	1	0
du	you	0	0	1	1
dr	doktor	0	0	1	0
dr	dr	0	0	1	0
dr	doctor	0	0	1	0
peyton	peyton	0	0	1	0
offret	the victim	0	0	1	0
offret	offering	0	0	1	0
runt	around	0	0	1	1
runt	between	0	0	1	0
emo	emo	0	0	1	0
humanism	humanistic	0	0	1	0
humanism	humanism	0	0	1	1
lärda	literate	0	0	1	0
lärda	scholars	0	0	1	0
lärda	savants	0	0	1	0
åka	go	0	0	1	1
åka	aka	0	0	1	0
helsingör	helsingor	0	0	1	0
helsingör	elsinore	0	0	1	0
helsingör	helsingör	0	0	1	0
sentida	recent	0	0	1	0
splittrades	shattered	0	0	1	0
splittrades	split	0	0	1	0
offren	victims	0	0	1	0
tyngre	heavy	0	0	1	0
tyngre	heavier	0	0	1	0
långhårig	rough	0	0	1	0
långhårig	long haired	0	0	1	0
långhårig	long-haired	0	0	1	1
utrotning	extinction	0	0	1	0
utrotning	extermination	0	0	1	1
libanon	lebanon	0	0	1	1
lärde	learned	0	0	1	0
kurdiska	kurdish	0	0	1	0
vanlig	ordinary	0	0	1	1
vanlig	common	0	0	1	1
vanlig	normal	0	0	1	0
treenigheten	tinity	0	0	1	0
treenigheten	the trinity	0	0	1	0
treenigheten	trinity	0	0	1	0
stewie	stewie	0	0	1	0
inne	inside	0	0	1	1
inne	in	0	0	1	1
avbryta	cancel	0	0	1	0
sexuell	sexual	0	0	1	1
djuret	the animal	0	0	1	0
djuret	animal	0	0	1	0
fornnordiska	old nordic	0	0	1	0
fornnordiska	ancient nordic	0	0	1	0
fornnordiska	old norse	0	0	1	0
piratpartiet	pirtpartiet	0	0	1	0
piratpartiet	pirate party	0	0	1	0
djuren	the animals	0	0	1	0
djuren	animals	0	0	1	0
materialet	the material	0	0	1	0
materialet	material	0	0	1	0
smaken	the flavour	0	0	1	0
smaken	flavor	0	0	1	0
osmanska	ottoman	0	0	1	0
osmanska	osmanian	0	0	1	0
osmanska	ottoman; osmanli	0	0	1	0
komplikationer	complications	0	0	1	0
we	we	0	0	1	0
intog	occupied	0	0	1	0
intog	seized	0	0	1	0
intog	took	0	0	1	0
dä	the elder	0	0	1	0
dä	with	0	0	1	0
då	then	0	0	1	1
då	when	0	0	1	1
dö	die	0	0	1	1
huvudsakligen	generally	0	0	1	0
huvudsakligen	primarily	0	0	1	0
försörjde	living	0	0	1	0
försörjde	provided	0	0	1	0
garanterar	ensures	0	0	1	0
garanterar	guarantees	0	0	1	0
muhammed	muhammed	0	0	1	0
cox	cox	0	0	1	1
gösta	gösta	0	0	1	0
gösta	gosta	0	0	1	0
medverkade	participated; contributed	0	0	1	0
medverkade	participated	0	0	1	0
kommer	is	0	0	1	0
fåfotingar	fÃ¥fotingar	1	0	1	0
fåfotingar	over	1	0	1	0
fåfotingar	pauropoda	1	1	0	0
fåfotingar	n/a	1	0	1	0
fåfotingar	arthropods	1	0	1	0
fåfotingar	dafotingar	1	0	1	0
fåfotingar	fafotingar	1	0	1	0
fåfotingar	centipede	1	0	1	0
fåfotingar	pauropods	1	0	1	0
väg	vague	0	0	1	0
väg	way	0	0	1	1
brad	brad	0	0	1	0
gruppens	group (-s)	0	0	1	0
gruppens	group	0	0	1	0
samverkan	co	0	0	1	0
samverkan	cooperation	0	0	1	1
graviditeten	the pregnacy	0	0	1	0
graviditeten	the pregnancy	0	0	1	0
väl	selecting	0	0	1	0
väl	good	0	0	1	0
vän	van	0	0	1	0
vän	friend	0	0	1	1
framgångsrikt	successful	0	0	1	0
framgångsrikt	successfully	0	0	1	1
någonting	nothing	0	0	1	0
någonting	anything	0	0	1	1
thierry	thierry	0	0	1	0
tusentals	thousands	0	0	1	0
framgångsrika	successful	0	0	1	0
framgångsrika	successes	0	0	1	0
framgångsrika	succesful	0	0	1	0
tony	tony	0	0	1	0
slaveriet	slavery	0	0	1	0
smith	smith	0	0	1	0
japans	japans	0	0	1	0
japans	japan's	0	0	1	0
patienten	patient	0	0	1	0
patienten	the patient	0	0	1	0
biologiska	biological	0	0	1	0
sjöar	lakes	0	0	1	0
sjöar	parks	0	0	1	0
begår	commits	0	0	1	0
begår	commit	0	0	1	0
hitlers	hitlers	0	0	1	0
patienter	patients	0	0	1	0
klubblag	club teams	0	0	1	0
klubblag	club team	0	0	1	0
spårvagnar	trams	0	0	1	0
spårvagnar	saving carriages	0	0	1	0
tillräckliga	insufficient	0	0	1	0
tillräckliga	sufficient	0	0	1	0
attacken	the attack	0	0	1	0
attacken	attack	0	0	1	0
fängelset	prison	0	0	1	0
fest	festival	0	0	1	1
fest	party	0	0	1	1
fest	fest	0	0	1	1
juridik	law	0	0	1	1
växthusgaser	vaxthusgaser	0	0	1	0
växthusgaser	greenhouse gas	0	0	1	0
drottningen	queen	0	0	1	0
drottningen	the queen	0	0	1	0
frekvens	frequencies	1	1	0	0
frekvens	freckvens	1	0	1	0
frekvens	value	1	0	1	0
frekvens	frequency	1	1	1	1
frekvens	date	1	0	1	0
frekvens	by number of	1	0	1	0
dödsstraffet	capital punishment; death penalty	0	0	1	0
dödsstraffet	death penalty	0	0	1	0
dödsstraffet	the death penalty	0	0	1	0
bulgariens	bulgaria	0	0	1	0
bulgariens	bulgaria's	0	0	1	0
fromstart	starting from	0	0	1	0
vagn	wagon	0	0	1	1
vagn	carrige	0	0	1	0
johansson	johansson	0	0	1	0
någonsin	ever	0	0	1	1
kupp	kupp	0	0	1	0
kupp	coup	0	0	1	1
kupp	coup (d'etat)	0	0	1	0
förändringarna	changes	0	0	1	0
förändringarna	change	0	0	1	0
aik	aik	0	0	1	0
tillväxten	growth	0	0	1	0
tillhandahåller	provides	0	0	1	0
klippa	cut	0	0	1	1
spanjorerna	spaniards	0	0	1	0
spanjorerna	spanish	0	0	1	0
spanjorerna	the spaniards	0	0	1	0
utanför	outside	0	0	1	1
vänt	turned	0	0	1	0
stålgemenskapen	steel community	0	0	1	0
minst	at least	0	0	1	0
lösa	solve	0	0	1	1
deltagarna	the participants	0	0	1	0
deltagarna	participants	0	0	1	0
frågade	inquired	0	0	1	0
frågade	asked	0	0	1	0
jordbruk	agricultural	0	0	1	0
tillträde	access	0	0	1	1
värderingar	evaluations	0	0	1	0
värderingar	values	0	0	1	0
löst	solved	0	0	1	1
löst	dissolved	0	0	1	0
löst	1st sentence: loosely; 2nd & 3rd: solved	0	0	1	0
rörelsen	movement	0	0	1	0
patent	patent	0	0	1	1
datorer	pc	0	0	1	0
bergskedjor	mountain ranges	0	0	1	0
föranledde	brought about	0	0	1	0
föranledde	led	0	0	1	0
utgår	deleted	0	0	1	0
utgivna	issued	0	0	1	0
utgivna	published	0	0	1	0
rörelser	movements	0	0	1	0
rörelser	movement	0	0	1	0
ersattes	was replaced by	0	0	1	0
ersattes	replaced	0	0	1	0
andelen	share	0	0	1	0
andelen	the share	0	0	1	0
andelen	the proportion	0	0	1	0
världsbanken	world bank	0	0	1	1
producerades	produced	0	0	1	0
producerades	was produced	0	0	1	0
platina	platinum	0	0	1	1
hann	did	0	0	1	0
hann	reached	0	0	1	0
hann	managed to (in a period of time)	0	0	1	0
saddam	saddam	0	0	1	0
balkan	balkan	0	0	1	0
balkan	the balkans	0	0	1	0
sexualitet	sexuality	0	0	1	1
delstater	states	0	0	1	0
hand	care	0	0	1	0
hand	hand	0	0	1	1
delstaten	land	0	0	1	0
delstaten	the state	0	0	1	0
hans	his	0	0	1	1
bilen	the car	0	0	1	0
bilen	car	0	0	1	0
koncentrerad	concentrated	0	0	1	1
koncentrerad	concentration	0	0	1	0
förföljelse	persecution	0	0	1	1
aspekter	aspects	0	0	1	0
sovjet	soviet	0	0	1	0
kyla	cold	0	0	1	1
kyla	cooling	0	0	1	0
riksdag	parliament; diet	0	0	1	0
riksdag	parliament	0	0	1	1
riksdag	the parliament	0	0	1	0
somliga	some people	0	0	1	0
somliga	some	0	0	1	1
styrkorna	forces	0	0	1	0
mamma	mother	0	0	1	1
monaco	monaco	0	0	1	0
dagar	says	0	0	1	0
dagar	day	0	0	1	0
dagar	days	0	0	1	0
the	the	0	0	1	0
thc	thc	0	0	1	0
skottland	scotland	0	0	1	1
använda	using	0	0	1	0
newton	newton	0	0	1	0
kall	cold	0	0	1	1
använde	used	0	0	1	0
bröder	brothers	0	0	1	0
kroppens	the body's	0	0	1	0
kroppens	the bodies	0	0	1	0
goda	good	0	0	1	0
enades	agreed	0	0	1	0
kalender	calendar	0	0	1	1
kalender	calender	0	0	1	0
swahili	swahili	0	0	1	0
swahili	swahilli	0	0	1	0
anställda	employed	0	0	1	0
distributioner	distributions	0	0	1	0
wright	wright	0	0	1	0
havets	the seas	0	0	1	0
havets	sea	0	0	1	0
skick	state	0	0	1	1
skick	condition	0	0	1	1
kvinnan	woman	0	0	1	0
kvinnan	female	0	0	1	0
plasma	plasma	0	0	1	1
viking	viking	0	0	1	1
maya	maya	0	0	1	0
rna	rna	0	0	1	0
skadorna	injuries	0	0	1	0
skadorna	damages	0	0	1	0
skadorna	damage	0	0	1	0
godkänna	approve	0	0	1	1
fusion	fusuion	0	0	1	0
fusion	fusion	0	0	1	1
indianer	indians	0	0	1	0
everton	everton	0	0	1	0
picasso	picasso	0	0	1	0
hepatit	hepatite	0	0	1	1
hepatit	hepatitis	0	0	1	1
hepatit	heptatitis	0	0	1	0
acceptera	acceptable	0	0	1	0
acceptera	accept	0	0	1	1
indelning	the subdivision	0	0	1	0
indelning	classification	0	0	1	0
indelningen	division	0	0	1	0
indelningen	subdivision	0	0	1	0
indelningen	classification	0	0	1	0
samfund	communities	0	0	1	0
samfund	order	0	0	1	0
°c	celsius	0	0	1	0
gandhi	gandhi	0	0	1	0
planeterna	the planet's	0	0	1	0
planeterna	planets	0	0	1	0
planeterna	the planets	0	0	1	0
transkription	transcription	0	0	1	1
transkription	transcript	0	0	1	0
transkription	transcripton	0	0	1	0
sixx	sixx	0	0	1	0
motsvarighet	equivalent	0	0	1	1
korea	koreans	0	0	1	0
korea	korea	0	0	1	1
utbröt	broke out	0	0	1	0
utbröt	erupted	0	0	1	0
populärkultur	popular culture	0	0	1	0
populärkultur	pop-culture	0	0	1	0
bort	away	0	0	1	1
bort	remove	0	0	1	0
färdiga	finished	0	0	1	0
färdiga	completed	0	0	1	0
born	born	0	0	1	0
presidentvalet	presidential elections	0	0	1	0
presidentvalet	presidential election	0	0	1	0
borg	tower	0	0	1	0
borg	castle	0	0	1	1
bord	table	0	0	1	1
händelser	handelsar	0	0	1	0
händelser	happenings	0	0	1	0
händelser	events	0	0	1	0
kungar	kings	0	0	1	0
humor	humor	0	0	1	1
humor	humour	0	0	1	1
territorierna	territories	0	0	1	0
purple	purple	0	0	1	0
sända	transmitting	0	0	1	0
sända	broadcast	0	0	1	0
sända	send	0	0	1	1
sände	sent	0	0	1	0
sände	limiting	0	0	1	0
rädd	scared	0	0	1	1
rädd	afraid	0	0	1	1
serbiens	serbias	0	0	1	0
siffran	the number	0	0	1	0
siffran	figure	0	0	1	0
siffran	number	0	0	1	0
sänds	sends	0	0	1	0
sänds	sands	0	0	1	0
sänds	sent	0	0	1	0
händelsen	the occurence	0	0	1	0
händelsen	event	0	0	1	0
vinterkriget	the winter war	0	0	1	0
vinterkriget	winter	0	0	1	0
vinterkriget	winter war	0	0	1	0
columbus	columbus	0	0	1	0
föredrar	prefer	0	0	1	0
föredrar	preferred	0	0	1	0
stadsdelarna	districts	0	0	1	0
stadsdelarna	neighborhood (-s)	0	0	1	0
skarsgård	skarsgård	0	0	1	0
skarsgård	cut farm	0	0	1	0
bevara	preserve	0	0	1	1
bevara	preserving	0	0	1	0
post	week	0	0	1	0
post	not a swedish word	0	0	1	0
detta	this	0	0	1	1
detta	that	0	0	1	0
detta	delta	0	0	1	0
vunnit	win	0	0	1	0
vunnit	won	0	0	1	0
innehållet	content	0	0	1	0
innehållet	contents	0	0	1	0
innehåller	contains	0	0	1	0
innehåller	include	0	0	1	0
införande	introduction	0	0	1	1
banker	banks	0	0	1	0
förhärskande	dominant	0	0	1	1
förhärskande	prevailing	0	0	1	0
olika	different	0	0	1	0
olika	variety	0	0	1	0
jacques	jacques	0	0	1	0
påstående	claim	0	0	1	0
påstående	assumption	0	0	1	0
påstående	pastilles of	0	0	1	0
samer	sami	0	0	1	0
istället	instead	0	0	1	0
istället	instead of	0	0	1	0
lois	lois	0	0	1	0
sedan	then	0	0	1	1
sedan	since	0	0	1	1
uppenbarelse	apparition	0	0	1	1
uppenbarelse	revelation	0	0	1	1
föddes	was born	0	0	1	0
föddes	born	0	0	1	0
blivande	prospective	0	0	1	1
blivande	future	0	0	1	1
blivande	to be	0	0	1	0
gemenskapen	the collective	0	0	1	0
gemenskapen	community	0	0	1	0
way	väg	0	0	1	0
way	way	0	0	1	0
dödsfall	death	0	0	1	1
dödsfall	deaths	0	0	1	0
was	was	0	0	1	0
war	war	0	0	1	0
beräknas	calculated	0	0	1	0
beräknas	estimated	0	0	1	0
beräknas	computed	0	0	1	0
expansionen	expansion	0	0	1	0
expansionen	the expansion	0	0	1	0
hypotes	hypothesized	0	0	1	0
hypotes	hypothesis	0	0	1	1
skiljas	separated	0	0	1	0
skiljas	separate	0	0	1	0
akondroplasi	archondroplasia	1	0	1	0
akondroplasi	created	1	0	1	0
akondroplasi	kondroplasia	1	1	0	0
akondroplasi	achodroplasia	1	0	1	0
akondroplasi	achondroplasia	1	1	0	0
akondroplasi	akondroplasia	1	1	0	0
förut	requires	0	0	1	0
förut	previously by	0	0	1	0
förut	before	0	0	1	1
moldavien	moldova	0	0	1	0
partiledare	party leader	0	0	1	0
ägnade	dedicated	0	0	1	0
ägnade	baited	0	0	1	0
emil	emil	0	0	1	0
reser	travels	0	0	1	0
reser	rise	0	0	1	0
reser	rises	0	0	1	0
studierna	studies	0	0	1	0
studierna	the studies	0	0	1	0
släppts	released	0	0	1	0
mtv	mtv	0	0	1	0
hästar	horses	0	0	1	0
närliggande	adjacent	0	0	1	0
närliggande	nearby	0	0	1	1
jämlikhet	equality	0	0	1	1
tvåa	second	0	0	1	1
väsen	being	0	0	1	1
väsen	vase	0	0	1	0
väsen	entity	0	0	1	1
engagerade	dedicated	0	0	1	0
engagerade	engaged	0	0	1	0
engagerade	committed	0	0	1	0
moore	moore	0	0	1	0
utomlands	abroad	0	0	1	1
tesla	tesla	0	0	1	0
xiis	xii	0	0	1	0
främmande	foreign; alien	0	0	1	0
främmande	undesirable	0	0	1	0
främmande	foreign	0	0	1	1
hölls	was held	0	0	1	0
hölls	was	0	0	1	0
efter	after	0	0	1	1
bilderna	the pictures	0	0	1	0
xiii	xiii	0	0	1	0
moln	cloud	0	0	1	1
moln	cloudy	0	0	1	0
empati	empathy	0	0	1	1
köket	cuisine	0	0	1	0
köket	the kitchen	0	0	1	0
blodtryck	blood pressure	0	0	1	1
toppen	top	0	0	1	0
toppen	peak	0	0	1	0
toppen	the top	0	0	1	0
alltid	always	0	0	1	1
arkitekten	architect	0	0	1	0
arkitekten	the architect	0	0	1	0
baháulláh	bahaullah	0	0	1	0
baháulláh	bahullah	0	0	1	0
järn	iron	0	0	1	1
järn	kon	0	0	1	0
arkitekter	architects	0	0	1	0
test	test	0	0	1	1
äger	owns	0	0	1	0
konservatism	conservatism	0	0	1	1
stränga	severe	0	0	1	0
femton	fifteen	0	0	1	1
tottenham	tottenham	0	0	1	0
reglerar	regulates	0	0	1	0
reglerar	controls	0	0	1	0
regleras	regulated	0	0	1	0
regleras	controlled	0	0	1	0
regleras	is regulated	0	0	1	0
definiera	defining	0	0	1	0
definiera	define	0	0	1	1
hemma	home	0	0	1	1
hemma	at home	0	0	1	1
omgivande	surrounding	0	0	1	0
omgivande	surounding	0	0	1	0
omgivande	ambient	0	0	1	1
solens	the sun	0	0	1	0
solens	solar	0	0	1	0
bergmans	bergman's	0	0	1	0
bergmans	bergmans	0	0	1	0
dance	dance	0	0	1	0
uppfanns	was invented	0	0	1	0
uppfanns	invented	0	0	1	0
tenderar	tend	0	0	1	0
datum	date	0	0	1	1
lider	suffering	0	0	1	0
lider	suffers	0	0	1	0
rättegången	trial	0	0	1	0
rättegången	the trial	0	0	1	0
rådde	prevailed	0	0	1	0
rådde	was	0	0	1	0
afrikaner	africans	0	0	1	0
släkting	relative	0	0	1	1
heller	neither	0	0	1	0
heller	neither; nor	0	0	1	0
heller	nor	0	0	1	0
igelkott	hedgehog	0	0	1	1
zone	zone	0	0	1	0
idén	the idea	0	0	1	0
idén	idea	0	0	1	0
terror	terror	0	0	1	0
tillstånd	state	0	0	1	1
tillstånd	to the dental	0	0	1	0
tillstånd	condition	0	0	1	1
hävdar	states	0	0	1	0
hävdar	assert	0	0	1	0
hävdar	maintain	0	0	1	0
hävdat	argued	0	0	1	0
hävdat	claimed	0	0	1	0
hannah	hannah	0	0	1	0
uttrycka	express	0	0	1	1
enskild	single	0	0	1	0
hannar	males	0	0	1	0
vegas	vegas	0	0	1	0
uttryckt	expressed	0	0	1	0
ölet	the beer	0	0	1	0
ölet	beer	0	0	1	0
enskilt	individually	0	0	1	0
enskilt	single	0	0	1	0
stycken	pieces; parts	0	0	1	0
stycken	pieces	0	0	1	0
gud	god	0	0	1	1
nedsatt	impaired	0	0	1	0
nedsatt	reduced	0	0	1	1
nedsatt	decreased; diminished	0	0	1	0
gul	yellow	0	0	1	1
levnadsstandard	living standard	0	0	1	0
levnadsstandard	standard of living	0	0	1	1
guy	guy	0	0	1	0
ljuset	the light	0	0	1	0
ljuset	light	0	0	1	0
formella	formal	0	0	1	0
templet	the temple	0	0	1	0
templet	temple	0	0	1	0
revolution	revolution	0	0	1	1
alfa	alpha	0	0	1	1
cosa	cosa	0	0	1	0
engagerad	dedicated	0	0	1	1
engagerad	engaged	0	0	1	1
invandrade	immigrated	0	0	1	0
invandrade	immigrant	0	0	1	0
väst	west	0	0	1	1
väst	the west	0	0	1	0
formellt	formally	0	0	1	1
formellt	formal	0	0	1	0
finländska	finish	0	0	1	0
finländska	finnish	0	0	1	0
motsatte	opposed	0	0	1	0
midsommar	midsummer	0	0	1	1
stimulera	stimulate	0	0	1	1
stimulera	stimulating	0	0	1	0
motsatta	opposite	0	0	1	0
yorks	yorks	0	0	1	0
ungdomar	youths	0	0	1	0
ungdomar	adolescents	0	0	1	0
ungdomar	the youth	0	0	1	0
tidig	early	0	0	1	1
ingick	were included	0	0	1	0
ingick	was	0	0	1	0
kosmiska	the cosmic	0	0	1	0
kosmiska	cosmic	0	0	1	0
uniform	uniform	0	0	1	1
fastigheter	real estates	0	0	1	0
fastigheter	properties	0	0	1	0
utspelar	takes place	0	0	1	0
utspelar	set	0	0	1	0
naturliga	natural	0	0	1	0
sökt	pending	0	0	1	0
sökt	searched	0	0	1	0
versionen	edition	0	0	1	0
versionen	the version	0	0	1	0
gener	genes	0	0	1	0
användbara	usable	0	0	1	0
användbara	useful	0	0	1	0
högst	highest	0	0	1	1
högst	maximum	0	0	1	0
marxismen	marxism	0	0	1	0
marxismen	the marxism	0	0	1	0
klassificeras	classified	0	0	1	0
klassificeras	lassificeras	0	0	1	0
genen	gene	0	0	1	0
genen	the gene	0	0	1	0
söka	search	0	0	1	1
söka	searching	0	0	1	0
människor	human	0	0	1	0
människor	people	0	0	1	0
näst	second	0	0	1	1
näst	second (to)	0	0	1	0
antarktiska	antarctic	0	0	1	0
flames	flames	0	0	1	0
kemi	chemistry	0	0	1	1
turné	tour	0	0	1	0
franklin	franklin	0	0	1	0
ponny	pony	0	0	1	1
fronten	front	0	0	1	0
fronten	the front	0	0	1	0
vinnare	win	0	0	1	0
vinnare	winner	0	0	1	1
ekr	ekr	0	0	1	0
ekr	ad	0	0	1	0
churchill	churchill	0	0	1	0
marken	soil	0	0	1	0
extra	optional	0	0	1	0
extra	extra	0	0	1	1
vapnet	the weapon	0	0	1	0
vapnet	the weapon; escutheon; coat of arms; arms; badge	0	0	1	0
spridit	spread	0	0	1	0
spridit	disseminated	0	0	1	0
ukrainas	ukranian	0	0	1	0
ukrainas	ukraine's	0	0	1	0
ukrainas	ukrainian	0	0	1	0
innebära	mean	0	0	1	0
vapnen	weapons	0	0	1	0
vapnen	the weapons	0	0	1	0
krigare	warriors	0	0	1	0
krigare	warrior	0	0	1	1
fbi	fbi	0	0	1	0
presenterar	presents	0	0	1	0
presenterar	present	0	0	1	0
presenteras	was presented	0	0	1	0
presenteras	presented	0	0	1	0
efterföljande	subsequent	0	0	1	0
territorier	territories	0	0	1	0
stabilitet	stability	0	0	1	1
live	live	0	0	1	1
regel	rule	0	0	1	1
motsvarar	comparable	0	0	1	0
motsvarar	corresponds to the	0	0	1	0
motsvarar	corresponds	0	0	1	0
angels	angels	0	0	1	0
parallellt	at the same time	0	0	1	0
parallellt	parallel	0	0	1	0
club	club	0	0	1	0
rivalitet	rivality	0	0	1	0
rivalitet	rivalry	0	0	1	1
snabbt	fast	0	0	1	1
snabbt	quickly	0	0	1	1
gärning	deed	0	0	1	1
gärning	enmeshing	0	0	1	0
motståndet	the resistance	0	0	1	0
motståndet	the resistence	0	0	1	0
parallella	parallel	0	0	1	0
zarathustra	zarathustra	0	0	1	0
västlig	western	0	0	1	0
länge	long	0	0	1	1
snabba	rapid	0	0	1	0
snabba	fast	0	0	1	0
användaren	the user	0	0	1	0
användaren	user	0	0	1	0
ibm	ibm	0	0	1	0
ibn	ibn	0	0	1	0
interaktion	the interaction	0	0	1	0
interaktion	interaction	0	0	1	1
frukt	fruit	0	0	1	1
frukt	fruits	0	0	1	0
can	can	0	0	1	0
can	cancer	0	0	1	0
erbjuder	offers	0	0	1	0
heart	heart	0	0	1	0
december	december	0	0	1	1
nobels	nobel's	0	0	1	0
nobels	nobel	0	0	1	0
influensavirus	flu virus	0	0	1	0
influensavirus	influenza	0	0	1	0
influensavirus	flue virus	0	0	1	0
gentemot	towards	0	0	1	1
gentemot	against	0	0	1	1
abort	abortion	0	0	1	1
ligan	league	0	0	1	0
pojke	boy	0	0	1	1
följas	followed	0	0	1	0
betydelse	importance	0	0	1	1
betydelse	eea	0	0	1	0
betydelse	significance	0	0	1	1
upprättades	was established	0	0	1	0
upprättades	establish	0	0	1	0
kopplingar	connections	0	0	1	0
kopplingar	links	0	0	1	0
perserna	the persians	0	0	1	0
perserna	persians	0	0	1	0
oändligt	infinity	0	0	1	0
oändligt	infinitely	0	0	1	0
southern	southern	0	0	1	0
kombattant	combatant	1	1	0	1
riktlinjer	guidelines	0	0	1	0
européerna	europeans	0	0	1	0
européerna	european	0	0	1	0
ungern	hungary	0	0	1	0
ungern	hungaria	0	0	1	0
stängt	closed	0	0	1	0
romarna	romans	0	0	1	0
romarna	the roman	0	0	1	0
romarna	the romans	0	0	1	0
flyttas	is moved	0	0	1	0
flyttas	moved	0	0	1	0
flyttar	move	0	0	1	0
värnplikt	military service	0	0	1	1
stänga	close	0	0	1	1
stänga	off	0	0	1	0
stänga	switch off	0	0	1	0
kurt	kurt	0	0	1	0
kurs	course	0	0	1	1
kurs	rate	0	0	1	1
michel	michel	0	0	1	0
ukrainska	ukrainian	0	0	1	0
rekordet	record	0	0	1	0
rekordet	the record	0	0	1	0
maktens	the powers	0	0	1	0
maktens	forces	0	0	1	0
maktens	the power's	0	0	1	0
ingripa	act	0	0	1	0
ingripa	interfere	0	0	1	1
ganska	rather	0	0	1	1
ganska	fairly	0	0	1	1
ganska	quite	0	0	1	1
grundades	founded	0	0	1	0
grundades	was founded	0	0	1	0
respektive	and	0	0	1	0
respektive	respective	0	0	1	1
mäter	measuring	0	0	1	0
mäter	measure	0	0	1	0
uppåt	raised	0	0	1	0
uppåt	up	0	0	1	1
uppåt	upwards	0	0	1	1
skabb	mites	0	0	1	0
skabb	scab	0	0	1	1
skabb	scabies	0	0	1	1
målningar	paintings	0	0	1	0
levde	lived	0	0	1	0
levde	survived	0	0	1	0
bergskedjan	mountain range	0	0	1	0
bergskedjan	the mountain group	0	0	1	0
nominerades	was nominated	0	0	1	0
nominerades	nominated	0	0	1	0
hals	throat	0	0	1	1
hals	neck	0	0	1	1
varav	of which	0	0	1	0
varav	which	0	0	1	0
arton	18	0	0	1	0
arton	eighteen	0	0	1	1
halv	half	0	0	1	1
biskop	bishop	0	0	1	1
nog	sufficiently	0	0	1	1
nog	enough	0	0	1	1
komponenter	components	0	0	1	0
terrorismen	terrorism	0	0	1	0
terrorismen	the terrorism	0	0	1	0
not	note	0	0	1	1
nou	nou	0	0	1	0
rakt	straight	0	0	1	1
now	now	0	0	1	0
hall	hall	0	0	1	1
frihet	freedom	0	0	1	1
james	james	0	0	1	0
antyder	indicates	0	0	1	0
svält	starvation	0	0	1	1
svält	starvations	0	0	1	0
stockholm	stockholm	0	0	1	0
stockholm	stocholm	0	0	1	0
januari	january	0	0	1	1
drog	draw	0	0	1	0
drog	pulled	0	0	1	1
drog	drug	0	0	1	1
aspergers	downs syndrome	0	0	1	0
aspergers	aspergers	0	0	1	0
em	em	0	0	1	0
em	european championship	0	0	1	0
el	el	0	0	1	0
en	a	0	0	1	1
citat	quote	0	0	1	1
ej	not	0	0	1	1
ej	no	0	0	1	0
ed	ed	0	0	1	0
eg	ec	0	0	1	0
utbrett	wide	0	0	1	0
utbrett	widespread	0	0	1	0
fördelning	distribution	0	0	1	1
ex	eg	0	0	1	0
ex	ex	0	0	1	0
känslan	feeling	0	0	1	0
känslan	the feeling	0	0	1	0
känslan	sense	0	0	1	0
eu	eu	0	0	1	0
et	et	0	0	1	0
resultera	result	0	0	1	0
fuglesang	fuglesang	0	0	1	0
tillämpar	administer	0	0	1	0
tillämpar	practice	0	0	1	0
tillämpar	administers	0	0	1	0
tillämpas	applied	0	0	1	0
er	you	0	0	1	1
er	your	0	0	1	1
album	album	0	0	1	1
teorier	theories	0	0	1	0
kortare	shorter	0	0	1	0
stallone	stallone	0	0	1	0
stånd	in the context: (make) the war happen	0	0	1	0
stånd	position	0	0	1	0
sevärdheter	attractions	0	0	1	0
koffein	caffeine	0	0	1	1
koffein	caffein	0	0	1	0
genetisk	genetic	0	0	1	1
författaren	the author	0	0	1	0
författaren	author	0	0	1	0
carl	carl	0	0	1	0
marina	marina	0	0	1	0
marina	marine	0	0	1	0
betraktades	considered	0	0	1	0
betraktades	regarded	0	0	1	0
myndigheterna	authorities	0	0	1	1
myndigheterna	the authorities	0	0	1	0
myndigheterna	the authoroties	0	0	1	0
british	british	0	0	1	0
jönköping	jönköping	0	0	1	0
jönköping	jonkoping	0	0	1	0
kategorisvenskspråkiga	category swedish-speaking	0	0	1	0
tillståndet	state	0	0	1	0
tillståndet	condition	0	0	1	0
tillståndet	the state	0	0	1	0
arbetsgivare	employers	0	0	1	0
blind	blind	0	0	1	1
blind	bank	0	0	1	0
blind	blank	0	0	1	0
xi	xi	0	0	1	0
hjälpt	helped	0	0	1	0
derivatan	derivative	0	0	1	0
derivatan	the derivative	0	0	1	0
fagocyt	fagocyt	1	0	1	0
fagocyt	fagocyte	1	0	1	0
fagocyt	phage	1	0	1	0
fagocyt	way	1	0	1	0
fagocyt	phagocyte	1	1	0	1
ring	ring	0	0	1	1
xv	xv	0	0	1	0
hjälpa	helping	0	0	1	0
bergqvist	bergqvist	0	0	1	0
omtvistat	disputed	0	0	1	0
omtvistat	contentious	0	0	1	0
omtvistat	controversial	0	0	1	0
konungarike	kingdom	0	0	1	1
desmond	desmond	0	0	1	0
svenske	swedish	0	0	1	0
sheen	sheen	0	0	1	0
dessutom	moreover	0	0	1	1
dessutom	furthermore	0	0	1	1
dessutom	additionally; likewise	0	0	1	0
dessutom	furthermore; moreover	0	0	1	0
satsningar	ventures	0	0	1	0
satsningar	investments	0	0	1	0
satsningar	resources	0	0	1	0
that	that	0	0	1	0
vattenkraft	water power	0	0	1	0
vattenkraft	hydro	0	0	1	0
vattenkraft	hydroelectric power	0	0	1	0
fascisterna	the fascists	0	0	1	0
fascisterna	the facists	0	0	1	0
fascisterna	fascists	0	0	1	0
than	than	0	0	1	0
television	television	0	0	1	1
europeisk	european	0	0	1	1
sidorna	the pages	0	0	1	0
sidorna	pages	0	0	1	0
utbyggda	expanded	0	0	1	0
utbyggda	expand	0	0	1	0
yttre	outer	0	0	1	1
primära	primary	0	0	1	0
träffade	met	0	0	1	0
grundad	founded	0	0	1	0
grundad	based	0	0	1	1
craig	craig	0	0	1	0
premier	premiums	0	0	1	0
statsminister	prime minister	0	0	1	1
faktor	factor	0	0	1	1
kairo	cairo	0	0	1	0
grundat	founded	0	0	1	0
grundat	(was) found	0	0	1	0
grundat	based	0	0	1	0
grundar	bases	0	0	1	0
grundar	based	0	0	1	0
grundas	is based	0	0	1	0
grundas	based	0	0	1	0
reologi	reologi	1	0	1	0
reologi	air	1	0	1	0
reologi	ether	1	0	1	0
reologi	reology	1	1	0	0
reologi	rheology	1	1	0	0
anger	indicates	0	0	1	0
anger	gives	0	0	1	0
slag	type	0	0	1	1
slag	kinds	0	0	1	0
fortsatte	continued	0	0	1	0
fortsatta	continued	0	0	1	0
förluster	loss	0	0	1	0
förluster	losses	0	0	1	0
etiopiska	ethiopian	0	0	1	0
etiopiska	etiopian	0	0	1	0
förlusten	loss; defeat	0	0	1	0
förlusten	loss	0	0	1	0
online	line	0	0	1	0
online	online	0	0	1	0
numera	now	0	0	1	0
numera	nowadays	0	0	1	1
santiago	santiago	0	0	1	0
successivt	successively	0	0	1	1
successivt	progressively	0	0	1	0
bekostnad	detriment	0	0	1	0
bekostnad	expense	0	0	1	1
america	america	0	0	1	0
michelle	michelle	0	0	1	0
nordöst	north east	0	0	1	0
nordöst	northeast	0	0	1	0
lyfter	lift	0	0	1	0
lyfter	lifts	0	0	1	0
lyfter	lifting	0	0	1	0
kampanil	phagocyte	1	0	1	0
kampanil	lock	1	0	1	0
kampanil	campanile	1	1	0	1
kampanil	kampanil	1	0	1	0
kampanil	bell tower	1	1	0	0
kampanil	castle	1	0	1	0
kampanil	bellfry; bell tower	1	1	0	0
berg	mountain(-s)	0	0	1	0
berg	mountain	0	0	1	1
nordligaste	northern	0	0	1	0
nordligaste	northermost	0	0	1	0
nordligaste	northernmost	0	0	1	0
parlamentets	the parliament's	0	0	1	0
parlamentets	parliament	0	0	1	0
jämte	next (to)	0	0	1	0
jämte	together with	0	0	1	1
jämte	plus	0	0	1	0
orsaka	cause	0	0	1	1
abraham	abraham	0	0	1	0
väska	kazan	1	0	1	0
väska	fluid	1	0	1	0
väska	bag	1	1	0	1
väska	leather case	1	1	0	0
väska	suitcase	1	0	1	0
väska	vasks	1	0	1	0
väska	its	1	0	1	0
väska	pan	1	0	1	0
skapats	was created	0	0	1	0
skapats	generated	0	0	1	0
doktor	doctor	0	0	1	1
doktor	phd	0	0	1	0
kyrkorna	churches	0	0	1	0
kyrkorna	the churches	0	0	1	0
trosbekännelsen	creed	0	0	1	0
trosbekännelsen	faith of confession	0	0	1	0
nazisternas	the nazi's	0	0	1	0
nazisternas	nazi	0	0	1	0
närmare	further	0	0	1	0
närmare	close to	0	0	1	0
marocko	morocco	0	0	1	0
marocko	marocco	0	0	1	0
rätter	dishes	0	0	1	0
rätten	right	0	0	1	0
rätten	the court	0	0	1	0
colombo	colombo	0	0	1	0
teori	theory	0	0	1	1
japansk	japansk	0	0	1	0
japansk	japanese	0	0	1	1
perfekt	perfect	0	0	1	1
mannens	man's	0	0	1	1
mannens	man	0	0	1	0
byggda	constructed	0	0	1	0
peang	clamp	1	0	1	0
peang	evolution	1	0	1	0
peang	forceps	1	0	1	0
peang	hemostatic clamp	1	0	1	0
peang	hemostatic forceps	1	0	1	0
peang	hemostat	1	1	0	0
peang	peang	1	0	1	0
förefaller	appear	0	0	1	0
förefaller	it seems	0	0	1	0
förefaller	appears	0	0	1	0
mästarna	the champions	0	0	1	0
mästarna	champions	0	0	1	0
mästarna	the masters	0	0	1	0
varmblod	warmblood	0	0	1	0
varmblod	warm-blooded	0	0	1	0
adolf	adolf	0	0	1	0
ansträngningar	effort	0	0	1	0
himmel	heaven	0	0	1	1
huskvarna	huskvarna	0	0	1	0
epoken	epoch	0	0	1	0
epoken	the epoch	0	0	1	0
dagbok	diary	0	0	1	1
dagbok	log	0	0	1	0
sierra	sierra	0	0	1	0
sydligaste	southernmost	0	0	1	0
sydligaste	most southern	0	0	1	0
tornet	tower	0	0	1	0
tornet	the tower	0	0	1	0
riddare	knight	0	0	1	1
samuel	samuel	0	0	1	1
självständigt	independent	0	0	1	0
självständigt	independently	0	0	1	1
självständigt	independant	0	0	1	0
ambitioner	ambitions	0	0	1	0
premiären	premiere	0	0	1	0
premiären	premier	0	0	1	0
marxistisk	marxist	0	0	1	0
marxistisk	marxistic	0	0	1	0
handlingar	actions	0	0	1	0
drabbas	affected	0	0	1	0
drabbas	suffer	0	0	1	0
drabbas	troubled with	0	0	1	0
facupen	fa cup	0	0	1	0
facupen	fa-cup	0	0	1	0
älgen	elk; moose	0	0	1	0
älgen	moose	0	0	1	0
älgen	alga	0	0	1	0
wembley	wembley	0	0	1	0
bushadministrationen	the bushadministration	0	0	1	0
bushadministrationen	the bush administration	0	0	1	0
bushadministrationen	bush administration	0	0	1	0
öresund	the sound	0	0	1	0
öresund	Øresund	0	0	1	0
slutet	end	0	0	1	0
osbourne	osbourne	0	0	1	0
lämnades	left	0	0	1	0
lämnades	was	0	0	1	0
lämnades	was lefted	0	0	1	0
väntan	awaiting	0	0	1	0
väntan	waiting	0	0	1	1
väntan	wait	0	0	1	1
stjärnor	stars	0	0	1	0
väntat	expected	0	0	1	0
väntas	expected	0	0	1	0
väntas	is expected	0	0	1	0
väntar	waiting	0	0	1	0
väntar	expect	0	0	1	0
sport	athletics	0	0	1	0
sport	sport	0	0	1	1
såsom	such as	0	0	1	0
såsom	like	0	0	1	1
katastrofer	disasters	0	0	1	0
katastrofer	catastrophes	0	0	1	0
depressionen	the depression	0	0	1	0
depressionen	depression	0	0	1	0
konstaterade	concluded	0	0	1	0
konstaterade	established	0	0	1	0
konstaterade	stated	0	0	1	0
populäraste	rated	0	0	1	0
populäraste	most popular	0	0	1	0
dödligt	lethal	0	0	1	0
dödligt	deadly	0	0	1	1
ladin	ladin	0	0	1	0
depressioner	recessions	0	0	1	0
depressioner	depressions	0	0	1	0
depressioner	depression	0	0	1	0
israels	israels	0	0	1	0
israels	israeli	0	0	1	0
israels	israel's	0	0	1	0
import	import	0	0	1	1
kommunismens	communism	0	0	1	0
kommunismens	the communisms	0	0	1	0
kommunismens	the communism's	0	0	1	0
katastrofen	catastrophy	0	0	1	0
katastrofen	the catastrophy	0	0	1	0
katastrofen	disaster	0	0	1	0
döttrar	daughters	0	0	1	0
yta	surface	0	0	1	1
dominerande	dominant	0	0	1	1
dominerande	dominating	0	0	1	1
dominerande	dominerande	0	0	1	0
ronja	ronja	0	0	1	0
personlighet	character	0	0	1	1
personlighet	personality	0	0	1	1
välfärd	wealth	0	0	1	0
välfärd	welfare	0	0	1	1
utgivningen	release	0	0	1	0
utgivningen	the publication	0	0	1	0
utgivningen	the release	0	0	1	0
verket	plant; indeed	0	0	1	0
verket	plant	0	0	1	0
verket	board	0	0	1	0
länkar	links	0	0	1	0
lånat	borrowed	0	0	1	0
verken	plants	0	0	1	0
verken	wroks	0	0	1	0
utgavs	was published	0	0	1	0
utgavs	published	0	0	1	0
comeback	comeback	0	0	1	1
folkräkning	census	0	0	1	1
folkräkning	head count	0	0	1	0
folkräkning	public shaving	0	0	1	0
förhållandevis	relatively	0	0	1	0
monicas	monica	0	0	1	0
monicas	monica's	0	0	1	0
popsångare	popsinger	0	0	1	0
popsångare	pop singer	0	0	1	0
representativ	representative	0	0	1	1
placerad	placed	0	0	1	1
placerad	disposed	0	0	1	0
handlar	is	0	0	1	0
handlar	concerns	0	0	1	0
kristinas	kristina's	0	0	1	0
kristinas	crisis thawed	0	0	1	0
propaganda	propaganda	0	0	1	1
feminismen	feminism	0	0	1	0
själen	soul	0	0	1	0
själen	the soul	0	0	1	0
nils	nils	0	0	1	0
comet	comet	0	0	1	0
låtarna	the songs	0	0	1	0
låtarna	songs	0	0	1	0
placerar	place	0	0	1	0
placerar	places	0	0	1	0
placeras	placed	0	0	1	0
järnvägar	failways	0	0	1	0
järnvägar	railways	0	0	1	0
järnvägar	rail	0	0	1	0
avskaffande	elimination	0	0	1	0
avskaffande	abolition	0	0	1	1
avskaffande	abolishment	0	0	1	1
regeringens	government	0	0	1	0
regeringens	government's	0	0	1	0
bomull	cotton	0	0	1	1
handlande	action	0	0	1	0
allmänt	generally	0	0	1	1
allmänt	generally; public	0	0	1	0
allmänt	commonly	0	0	1	1
oliver	olives	0	0	1	0
lyssnade	listened	0	0	1	0
karlstads	karlstad's	0	0	1	0
sker	happens	0	0	1	0
sker	is	0	0	1	0
oden	node	0	0	1	0
oden	oden	0	0	1	0
knappt	barely	0	0	1	0
petit	petit	0	0	1	0
djurgården	djurgården	0	0	1	0
djurgården	zoo	0	0	1	0
ändrade	changed	0	0	1	0
ändrade	modified	0	0	1	0
krona	crown	0	0	1	1
observera	note	0	0	1	1
observera	observe	0	0	1	1
riktningar	directions	0	0	1	0
riktningar	direction	0	0	1	0
riktningar	direction (-s)	0	0	1	0
elvis	elvis	0	0	1	0
funnits	found	0	0	1	0
funnits	been	0	0	1	0
lösningsmedel	solvent	0	0	1	1
empathy	empathy	0	0	1	0
förbud	ban	0	0	1	1
förbud	prohibiting	0	0	1	0
förbud	prohibition	0	0	1	1
ytan	the area	0	0	1	0
ytan	surface	0	0	1	0
ytan	area	0	0	1	0
uefacupen	the uefa champions league	0	0	1	0
uefacupen	uefa europa league	0	0	1	0
uefacupen	uefacupen	0	0	1	0
ändringar	edit	0	0	1	0
ändringar	starts to process	0	0	1	0
ändringar	changes	0	0	1	0
prinsessan	the princess	0	0	1	0
prinsessan	princess	0	0	1	0
rapporten	report	0	0	1	0
rapporten	the report	0	0	1	0
polens	polands	0	0	1	0
polens	pole	0	0	1	0
ordningen	the order	0	0	1	0
ordningen	order	0	0	1	0
ordningen	procedure	0	0	1	0
motorvägarna	highways	0	0	1	0
motorvägarna	the highways	0	0	1	0
ansikte	face	0	0	1	1
tjeckien	czech republic	0	0	1	0
tjeckien	the czech republic	0	0	1	0
utfört	done	0	0	1	0
utförs	is done	0	0	1	0
utförs	out	0	0	1	0
föll	fell	0	0	1	0
förlängningen	elongation	0	0	1	0
förlängningen	forlajgningen	0	0	1	0
inslag	impact	0	0	1	0
inslag	elements	0	0	1	0
inslag	element	0	0	1	1
finanskrisen	financial crisis	0	0	1	0
finanskrisen	the financial crisis	0	0	1	0
behandlade	was treated	0	0	1	0
behandlade	treated	0	0	1	0
utförd	completed	0	0	1	0
utförd	performed	0	0	1	0
utföra	perform	0	0	1	1
utföra	out	0	0	1	0
kvarter	quarter	0	0	1	1
kvarter	neighborhoods	0	0	1	0
kvarter	block	0	0	1	1
kenya	kenya	0	0	1	1
katalanska	catalan	0	0	1	0
helium	helium	0	0	1	1
grundade	founded	0	0	1	0
grundade	based	0	0	1	0
slaget	the strike	0	0	1	0
slaget	type	0	0	1	0
orsakade	caused	0	0	1	0
orsakade	causing	0	0	1	0
programvara	software	0	0	1	1
självständighet	independance	0	0	1	0
självständighet	independence	0	0	1	1
media	media	0	0	1	1
iväg	away	0	0	1	0
iväg	off	0	0	1	0
misstänkt	accused	0	0	1	0
misstänkt	suspect	0	0	1	1
misstänkt	suspected of	0	0	1	0
talmannen	president	0	0	1	0
talmannen	speaker of the riksdag	0	0	1	0
homosexualitet	homosexuality	0	0	1	1
homosexualitet	homosexuallity	0	0	1	0
kromosom	chromosome	0	0	1	1
pesten	death	0	0	1	0
pesten	the plague	0	0	1	0
pesten	plague	0	0	1	0
lite	little	0	0	1	0
lite	a little	0	0	1	0
utför	perform	0	0	1	0
utför	out	0	0	1	0
figurer	figures	0	0	1	0
speciella	special	0	0	1	0
offensiven	offensive	0	0	1	0
offensiven	the offensive	0	0	1	0
ägdes	owned	0	0	1	0
skivbolaget	record label	0	0	1	0
skivbolaget	the record company	0	0	1	0
acdc	ac/dc	0	0	1	0
omfattande	wide-ranging	0	0	1	0
omfattande	large	0	0	1	1
omfattande	massive; extensive	0	0	1	0
omfattar	encompass	0	0	1	0
omfattar	include	0	0	1	0
omfattas	comprise	0	0	1	0
omfattas	subject	0	0	1	0
speciellt	particularly	0	0	1	1
speciellt	sppeciellt	0	0	1	0
förutsättningarna	prerequisites	0	0	1	0
förutsättningarna	conditions	0	0	1	0
ekonomisk	economic	0	0	1	1
tradition	tradition	0	0	1	1
undersökning	study	0	0	1	0
undersökning	survey	0	0	1	1
fredspris	peace prize	0	0	1	1
överhöghet	supremacy	0	0	1	1
överhöghet	suzeranity	0	0	1	0
överhöghet	sovereignty	0	0	1	0
in	in the context: recorded = spela (in)	0	0	1	0
in	in	0	0	1	1
stämmer	(if it's) true	0	0	1	0
stämmer	correct	0	0	1	0
stämmer	is true	0	0	1	0
användandet	usage	0	0	1	0
användandet	use	0	0	1	0
sträcka	distance	0	0	1	1
flaggor	flags	0	0	1	0
låga	cook	0	0	1	0
låga	low	0	0	1	0
mynning	outfall	0	0	1	1
mynning	muzzle	0	0	1	1
mynning	mouth	0	0	1	1
forskarna	the scientists	0	0	1	0
forskarna	scientists	0	0	1	0
skandinaviska	scandinavic	0	0	1	0
skandinaviska	scandinavian	0	0	1	0
tydlig	clear	0	0	1	1
tydlig	obvious	0	0	1	1
petter	petter	0	0	1	0
samiska	sami	0	0	1	0
eleverna	the pupils	0	0	1	0
eleverna	the students	0	0	1	0
allmänhet	in general	0	0	1	0
allmänhet	public	0	0	1	1
allmänhet	general	0	0	1	0
lagerkvist	lagerkvist	0	0	1	0
nazismen	nazism	0	0	1	0
euron	the euro	0	0	1	0
euron	euro	0	0	1	0
ca	cirka	0	0	1	0
ca	approximately	0	0	1	0
lade	laid	0	0	1	0
lade	added	0	0	1	0
lade	seized	0	0	1	0
ditt	your	0	0	1	0
irland	irland	0	0	1	0
irland	ireland	0	0	1	1
arbeta	work	0	0	1	1
arbeta	working	0	0	1	0
härifrån	from here	0	0	1	0
härifrån	here	0	0	1	0
stund	while	0	0	1	1
stund	momentum	0	0	1	0
selma	selma	0	0	1	0
amy	amy	0	0	1	0
medförde	resulted	0	0	1	0
medförde	brought	0	0	1	0
medförde	led	0	0	1	0
lady	lady	0	0	1	1
tobak	tobacco	0	0	1	1
nationella	national	0	0	1	0
skilda	seperated	0	0	1	0
skilda	separate	0	0	1	0
miniatyr|en	thumbnail	0	0	1	0
miniatyr|en	a minature	0	0	1	0
skilde	divided	0	0	1	0
skilde	varied	0	0	1	0
skilde	there was a separation	0	0	1	0
direktör	director	0	0	1	1
varandra	each other	0	0	1	1
nationellt	national	0	0	1	0
nationellt	nationally	0	0	1	0
t	t	0	0	1	0
t	e.g.	0	0	1	0
löner	wages and salaries	0	0	1	0
löner	salaries	0	0	1	0
astronomer	astronomers	0	0	1	0
astronomer	astronomer	0	0	1	0
inriktade	oriented	0	0	1	0
pjäs	piece	0	0	1	1
kategoripersoner	category of persons	0	0	1	0
berodde	was	0	0	1	0
berodde	depended	0	0	1	0
berodde	depended upon	0	0	1	0
säsongens	season	0	0	1	0
säsongens	the seasons	0	0	1	0
fråga	ask	0	0	1	1
fråga	fraga	0	0	1	0
fråga	question	0	0	1	1
agera	act	0	0	1	1
utskott	organ	0	0	1	0
utskott	committee	0	0	1	1
nsdap	nsdap	0	0	1	0
inuti	inside	0	0	1	1
kaffet	coffee	0	0	1	0
kaffet	the coffee	0	0	1	0
francis	francis	0	0	1	0
drama	drama	0	0	1	1
ideologi	ideology	0	0	1	1
läget	position	0	0	1	0
läget	location	0	0	1	0
central	central	0	0	1	1
central	center	0	0	1	1
nordliga	northernly	0	0	1	0
nordliga	northern	0	0	1	0
läger	camps	0	0	1	0
läger	camp	0	0	1	1
sri	sri	0	0	1	0
torget	square	0	0	1	0
torget	the square	0	0	1	0
torget	torget	0	0	1	0
bidragen	the contributions	0	0	1	0
bidragen	contributions	0	0	1	0
övergav	abandoned	0	0	1	0
efterkrigstiden	the post-war period	0	0	1	0
efterkrigstiden	post-war era	0	0	1	0
efterkrigstiden	post-war	0	0	1	0
söndagen	sunday	0	0	1	0
kapten	captain	0	0	1	1
klassiker	classics	0	0	1	0
klassiker	classic	0	0	1	1
transporter	carriage	0	0	1	0
transporter	transports	0	0	1	0
lissabonfördraget	treaty of lisbon	0	0	1	0
lissabonfördraget	lisbon treaty	0	0	1	0
your	your	0	0	1	0
fast	solid	0	0	1	1
fast	even though	0	0	1	0
fast	though; although; fixed; permanent	0	0	1	0
area	area	0	0	1	1
satsade	invested	0	0	1	0
satsade	bet	0	0	1	0
specifikt	specifically	0	0	1	0
stark	strong	0	0	1	1
dödade	killed	0	0	1	0
specifika	specific	0	0	1	0
småland	smaland	0	0	1	0
småland	småland	0	0	1	0
hawking	hawking	0	0	1	0
därför	because	0	0	1	0
därför	therefore	0	0	1	1
tillväxt	growth	0	0	1	1
wailers	wailers	0	0	1	0
infördes	introduced	0	0	1	0
infördes	were implemented	0	0	1	0
hälft	half	0	0	1	1
införde	enforced	0	0	1	0
införde	introduced	0	0	1	0
expeditionen	the expidition	0	0	1	0
expeditionen	expedition	0	0	1	0
minne	memory	0	0	1	1
engelskan	the english	0	0	1	0
engelskan	english	0	0	1	0
sålunda	thus	0	0	1	1
indelningar	divisions	0	0	1	0
indelningar	classifications	0	0	1	0
freddy	freddy	0	0	1	0
förbundsrepubliken	the federal republic	0	0	1	0
förbundsrepubliken	federal republic of	0	0	1	0
förbundsrepubliken	federal republic	0	0	1	0
miguel	miguel	0	0	1	0
expeditioner	expeditions	0	0	1	0
kostar	costs	0	0	1	0
kungen	king	0	0	1	0
kungen	the king	0	0	1	0
grammis	grammy	0	0	1	0
sveriges	swedens	0	0	1	0
sveriges	sweden	0	0	1	0
styrde	steered	0	0	1	0
knut	knut	0	0	1	0
knut	knot	0	0	1	1
transportera	transport	0	0	1	1
nere	down	0	0	1	1
nere	low	0	0	1	1
antropogen	conference	1	0	1	0
antropogen	ntropogen	1	0	1	0
antropogen	antropog	1	1	0	0
antropogen	an anthropogenic	1	1	0	0
antropogen	anthropogeny	1	0	1	0
antropogen	antropogenic	1	1	0	0
antropogen	created by humans	1	1	0	0
antropogen	man-made	1	0	1	0
antropogen	anthropogenic	1	1	0	0
drycker	beverages	0	0	1	0
mäktiga	powerful	0	0	1	0
självstyrande	self-governing	0	0	1	1
självstyrande	independent	0	0	1	0
självstyrande	self-governance	0	0	1	0
fortsätter	continues	0	0	1	0
fortsätter	continue	0	0	1	0
upphovsman	author	0	0	1	1
upphovsman	creator	0	0	1	1
you	you	0	0	1	0
mörker	dark	0	0	1	1
mörker	darkness	0	0	1	1
malmös	malmö	0	0	1	0
malmös	malmö's	0	0	1	0
bestående	comprising	0	0	1	0
bestående	lasting	0	0	1	1
drift	operation	0	0	1	1
drift	drift	0	0	1	1
bidragande	contributors	0	0	1	0
massachusetts	massachusetts	0	0	1	1
massachusetts	massachussetts	0	0	1	0
bandmedlemmarna	band members	0	0	1	0
bandmedlemmarna	have	0	0	1	0
anläggningar	plants	0	0	1	0
anläggningar	facilities	0	0	1	0
skuggan	shadow	0	0	1	0
skuggan	the shadow	0	0	1	0
mänsklighetens	humanity's	0	0	1	0
mänsklighetens	humanities	0	0	1	0
intåg	entry	0	0	1	1
intåg	advent	0	0	1	0
morgonen	the morning	0	0	1	0
morgonen	am	0	0	1	0
kläder	clades	0	0	1	0
kläder	clothes	0	0	1	1
föremål	object	0	0	1	1
föremål	subject	0	0	1	1
skådespelerska	actress	0	0	1	1
export	export	0	0	1	1
olympiastadion	olympa stadium	0	0	1	0
olympiastadion	olympic stadium	0	0	1	0
monte	assembly	0	0	1	0
eriksson	eriksson	0	0	1	0
beskrivningar	description	0	0	1	0
beskrivningar	descriptions	0	0	1	0
läste	read	0	0	1	0
messi	messi	0	0	1	0
loppet	bore	0	0	1	0
loppet	the race	0	0	1	0
atlanta	atlanta	0	0	1	0
antoinette	antoinette	0	0	1	0
hävda	claim	0	0	1	1
hävda	asserting	0	0	1	0
där	where	0	0	1	1
där	in which	0	0	1	0
där	were	0	0	1	0
foster	embryo	1	1	0	0
foster	mrs. foster	1	0	1	0
foster	infant	1	0	1	0
foster	fetus	1	1	1	1
foster	fetuses	1	0	1	0
foster	foster	1	0	1	0
foster	do not need	1	0	1	0
foster	nothing	1	0	1	0
foster	fomentar	1	0	1	0
foster	embryonic	1	0	1	0
foster	fetal	1	0	1	0
nästa	next	0	0	1	1
klorofyll	chlorophyll	0	0	1	1
klorofyll	cholophyll	0	0	1	0
vers	verse	0	0	1	1
jensen	jensen	0	0	1	0
vägrar	refuses	0	0	1	0
vägrar	refuse	0	0	1	0
kvinna	woman	0	0	1	1
ändrat	changed	0	0	1	0
ändrat	modified	0	0	1	0
verk	work	0	0	1	1
verk	works	0	0	1	0
osv	etc.	0	0	1	0
uppfattar	sees	0	0	1	0
uppfattar	percieves	0	0	1	0
uppfattar	interpret	0	0	1	0
tredje	third	0	0	1	1
heaven	heaven	0	0	1	0
sverige	sweden	0	0	1	1
louis	louis	0	0	1	0
tvskådespelare	tv actor	0	0	1	0
manager	manager	0	0	1	0
industrialiseringen	indutrialization	0	0	1	0
industrialiseringen	industrialization	0	0	1	0
tigern	tiger	0	0	1	0
tigern	the tiger	0	0	1	0
resan	the trip	0	0	1	0
resan	journey	0	0	1	0
uppfattas	be perceived	0	0	1	0
uppfattas	perceived	0	0	1	0
uppfattas	are regarded	0	0	1	0
rasism	racism	0	0	1	1
magdalena	magdalena	0	0	1	0
uppfylla	satisfy	0	0	1	1
uppfylla	fulfill	0	0	1	1
uppfylla	meet (requirements)	0	0	1	0
skiva	record	0	0	1	1
skiva	disc	0	0	1	1
egendom	property	0	0	1	1
kritiserats	criticized	0	0	1	0
kritiserats	critized	0	0	1	0
orgasm	orgasm	0	0	1	1
markerade	selected	0	0	1	0
markerade	marked	0	0	1	0
trupper	troops	0	0	1	0
bedrev	conducted	0	0	1	0
bedrev	managed	0	0	1	0
känna	known	0	0	1	0
känna	know	0	0	1	1
hår	hair	0	0	1	1
flög	fly	0	0	1	0
flög	flew	0	0	1	0
känns	feels	0	0	1	0
känns	felt	0	0	1	0
känns	feels like	0	0	1	0
föreställande	depicting	0	0	1	0
bernhard	bernhard	0	0	1	0
hål	hole	0	0	1	1
hål	hal	0	0	1	0
sattes	was added	0	0	1	0
inblandad	mixed	0	0	1	0
irak	iraq	0	0	1	1
ersatt	replaced	0	0	1	0
iran	iran	0	0	1	1
händer	happens	0	0	1	1
händer	happening	0	0	1	0
händer	hands	0	0	1	0
hålet	hole; gap	0	0	1	0
hålet	hole	0	0	1	0
hålet	the hole	0	0	1	0
kronor	kronor	0	0	1	0
kronor	crowns	0	0	1	0
observeras	observed	0	0	1	0
observeras	is noticed	0	0	1	0
observeras	is observed	0	0	1	0
uttalat	pronounced	0	0	1	0
uttalat	outspoken	0	0	1	0
uttalat	expressed	0	0	1	0
uttalas	pronounced	0	0	1	0
uttalas	be pronounced	0	0	1	0
arena	arena	0	0	1	1
medarbetare	employees	0	0	1	0
medarbetare	coworker	0	0	1	0
tillsätts	added	0	0	1	0
tillsätts	appointed	0	0	1	0
tillsätts	appoints	0	0	1	0
signifikant	significant	0	0	1	1
krigen	the wars	0	0	1	0
krigen	wars	0	0	1	0
dyker	dives	0	0	1	0
dyker	shows	0	0	1	0
renässansen	the renaissance	0	0	1	0
renässansen	renaissance	0	0	1	0
härkomst	origin	0	0	1	1
härkomst	provenance	0	0	1	0
boxning	boxing	0	0	1	1
boxning	boxing; pugilism	0	0	1	0
sagor	fairytales	0	0	1	0
sagor	tales	0	0	1	0
sagor	fairy tales	0	0	1	0
kriget	the war	0	0	1	0
kriget	war	0	0	1	0
hoppades	hoped	0	0	1	1
perspektiv	perspective	0	0	1	1
medicin	medicine	0	0	1	1
globen	lobe	0	0	1	0
globen	the globe	0	0	1	0
nazityskland	nazi germany	0	0	1	0
läst	read	0	0	1	0
läst	load	0	0	1	0
gick	went	0	0	1	0
gick	passed	0	0	1	0
grunda	found	0	0	1	1
grunda	base	0	0	1	1
dalarna	valleys	0	0	1	0
dalarna	dalarna	0	0	1	0
nukleotider	nucleotides	0	0	1	0
nukleotider	nucleotide	0	0	1	0
familj	family	0	0	1	1
avsedd	adapted	0	0	1	0
avsedd	intended	0	0	1	1
nathan	nathan	0	0	1	0
simba	simba	0	0	1	0
simba	pool	0	0	1	0
läsa	read	0	0	1	1
arrangemang	arrangement	0	0	1	1
taket	the roof	0	0	1	0
taket	ceiling	0	0	1	0
etablerad	established	0	0	1	1
spindlingar	slindlingar	1	0	1	0
spindlingar	fungal genus	1	1	0	0
spindlingar	cortinariuses	1	0	1	0
spindlingar	webcap	1	0	1	0
spindlingar	spindlingar	1	0	1	0
spindlingar	fungus	1	0	1	0
spindlingar	stalin	1	0	1	0
spindlingar	cortinarus	1	0	1	0
spindlingar	spiders	1	0	1	0
spindlingar	cortinarius	1	1	0	0
spindlingar	cortinariaceae	1	1	0	0
spindlingar	this is not a swedish word.	1	0	1	0
trummisen	the drummer	0	0	1	0
trummisen	drummer	0	0	1	0
oecd	oecd	0	0	1	0
bolagets	company's	0	0	1	0
bolagets	the corporation's	0	0	1	0
bolagets	company	0	0	1	0
representeras	represented	0	0	1	0
representerar	represents	0	0	1	0
förvaras	stored	0	0	1	0
förvaras	is stored	0	0	1	0
förvaras	material is kept	0	0	1	0
teatrar	theaters	0	0	1	0
massan	mass	0	0	1	0
kurdistan	kurdistan	0	0	1	0
tillbehör	sides	0	0	1	0
tillbehör	condiments	0	0	1	0
tillbehör	accessory	0	0	1	0
säljas	is sold	0	0	1	0
säljas	sold	0	0	1	0
kärleken	love	0	0	1	0
kärleken	find love	0	0	1	0
kärleken	the love	0	0	1	0
latinamerikanska	latin-american	0	0	1	0
latinamerikanska	latin american	0	0	1	0
längtan	longing	0	0	1	1
vm	world championship	0	0	1	0
vm	vm	0	0	1	0
inspelad	recorded	0	0	1	1
få	have; make; few	0	0	1	0
få	gain	0	0	1	1
få	fa	0	0	1	0
laryngoskop	evolution	1	0	1	0
laryngoskop	laryngoscope	1	1	0	1
laryngoskop	laryngoscopy	1	1	0	0
laryngoskop	llaryngoscope	1	0	1	0
laryngoskop	laryngoscopes	1	0	1	0
laryngoskop	laryngoskop	1	1	0	0
lagstiftande	legislative	0	0	1	1
lagstiftande	legislating	0	0	1	0
lagstiftande	legislation	0	0	1	0
nina	nina	0	0	1	0
gazaremsan	gaza strip	0	0	1	0
gazaremsan	the gaza strip	0	0	1	0
ombord	onboard	0	0	1	1
ombord	board	0	0	1	0
history	history	0	0	1	0
rapporterade	reported	0	0	1	0
feministiska	feminist	0	0	1	0
partner	partner	0	0	1	1
herrens	lord	0	0	1	0
species	species	0	0	1	0
zanzibar	zanzibar	0	0	1	0
serber	serbs	0	0	1	0
ledger	ledger	0	0	1	0
smitta	infection	0	0	1	1
reidars	reidars	0	0	1	0
reidars	reidar's	0	0	1	0
ytterligare	further	0	0	1	1
ytterligare	additional	0	0	1	1
samarbetet	co	0	0	1	0
samarbetet	cooperation	0	0	1	0
samarbetet	the collaboration	0	0	1	0
hustrun	the wife	0	0	1	0
hustrun	his wife	0	0	1	0
turkarna	turks	0	0	1	0
turkarna	the turks	0	0	1	0
torde	could	0	0	1	0
torde	should	0	0	1	1
maffia	mob	1	1	0	0
maffia	mafia	1	1	0	0
maffia	the mob	1	0	1	0
maffia	clinically	1	0	1	0
maffia	clinical	1	0	1	0
fc	fc	0	0	1	0
fd	former	0	0	1	0
fd	ex	0	0	1	0
ff	ff	0	0	1	0
invasion	invasions	0	0	1	0
invasion	invasion	0	0	1	1
samarbeten	cooperations	0	0	1	0
samarbeten	collaborations	0	0	1	0
fn	un	0	0	1	0
fn	the un	0	0	1	0
fn	fn	0	0	1	0
stabil	stable	0	0	1	1
däremot	on the contrary	0	0	1	1
däremot	however	0	0	1	0
västvärlden	west	0	0	1	0
västvärlden	western world	0	0	1	0
kostnaden	cost	0	0	1	0
byggandet	construction	0	0	1	0
byggandet	the building	0	0	1	0
skivan	record	0	0	1	0
skivan	the record	0	0	1	0
skivan	disc	0	0	1	0
enzymer	enzymes	0	0	1	0
korset	cross	0	0	1	0
vågen	the wave	0	0	1	0
vågen	scale	0	0	1	0
kognitiv	cognitive	0	0	1	1
segrar	wins	0	0	1	0
segrar	victories	0	0	1	0
kategoriorter	category visited	0	0	1	0
ö	island	0	0	1	1
ö	o	0	0	1	0
kostnader	cost	0	0	1	0
kostnader	costs	0	0	1	1
kostnader	expenses	0	0	1	0
dream	dream	0	0	1	0
släpps	released	0	0	1	0
släpps	(is) released	0	0	1	0
helt	completely	0	0	1	1
helt	totally	0	0	1	0
förlorades	lost	0	0	1	0
förlorades	was lost	0	0	1	0
bloggar	blogs	0	0	1	0
gångna	past	0	0	1	0
gångna	past; gone	0	0	1	0
helgdagar	holidays	0	0	1	0
tornen	towers	0	0	1	0
tornen	the tower	0	0	1	0
hela	entire	0	0	1	0
hela	full	0	0	1	0
maffian	mafia	0	0	1	0
hell	hell	0	0	1	0
kombinerade	combined	0	0	1	0
eros	eros	0	0	1	0
hundratusentals	hundreds of thousands of	0	0	1	0
hundratusentals	hundreds of thousands	0	0	1	1
paulo	paulo	0	0	1	0
hendrix	hendrix	0	0	1	0
antagits	adoption	0	0	1	0
antagits	adopted	0	0	1	0
systems	systems	0	0	1	0
systems	system	0	0	1	0
mahatma	mahatma	0	0	1	0
musikalisk	musical	0	0	1	1
bytte	changed	0	0	1	0
bytte	changed it's	0	0	1	0
bytte	swapped	0	0	1	0
trycket	pressure	0	0	1	0
konstitutionella	constitutional	0	0	1	0
greps	was arrested	0	0	1	0
greps	arrested	0	0	1	0
greps	(was) arrested	0	0	1	0
dyrt	a high price	0	0	1	0
dyrt	expensive	0	0	1	1
dyrt	dearly	0	0	1	1
västliga	western	0	0	1	0
fullt	full; fully; completely	0	0	1	0
fullt	completely	0	0	1	1
fullt	full	0	0	1	1
riksrådet	privy council	0	0	1	0
riksrådet	privy council; council of state; crown council; senate	0	0	1	0
riksrådet	riskradet	0	0	1	0
skådespelaren	actor	0	0	1	0
fulla	full	0	0	1	0
fulla	complete	0	0	1	0
förbättra	improve	0	0	1	1
skrivit	written	0	0	1	0
skrivit	wrote	0	0	1	0
die	die	0	0	1	0
kontinentens	the continents	0	0	1	0
kontinentens	continent	0	0	1	0
frånträde	relinquishment	0	0	1	0
frånträde	withdrawal	0	0	1	0
ifk	ifk	0	0	1	0
etnisk	ethnic	0	0	1	1
statyn	the statue	0	0	1	0
statyn	statue	0	0	1	0
neil	neil	0	0	1	0
positionen	position	0	0	1	0
positionen	the position	0	0	1	0
säljande	selling	0	0	1	1
äldste	elders	0	0	1	0
äldste	eldest	0	0	1	0
positioner	positions	0	0	1	0
låta	let	0	0	1	1
ersätts	replaced	0	0	1	0
överlägset	far	0	0	1	0
överlägset	superior	0	0	1	0
robert	robert	0	0	1	0
bodde	lived	0	0	1	0
ersätta	replacing	0	0	1	0
ersätta	replace	0	0	1	1
tilläts	was allowed	0	0	1	0
tilläts	were allowed to	0	0	1	0
tilläts	allowed	0	0	1	0
lungorna	lungs	0	0	1	0
lungorna	the lungs	0	0	1	0
pythagoras	pythagoras	0	0	1	0
återigen	once again	0	0	1	0
återigen	yet again	0	0	1	0
återigen	aterigen	0	0	1	0
utredningen	investigation	0	0	1	0
utredningen	the investigation	0	0	1	0
heroin	heroin	0	0	1	1
heroin	heroine	0	0	1	0
skönhet	beauty	0	0	1	1
delningen	division	0	0	1	0
delningen	pitch	0	0	1	0
vasas	vasa	0	0	1	0
vasas	vasas	0	0	1	0
vasas	vasa's	0	0	1	0
svarade	answered	0	0	1	0
svarade	said	0	0	1	0
svarade	accounted (for); answered	0	0	1	0
spets	edge; top	0	0	1	0
spets	tip	0	0	1	1
spets	point	0	0	1	1
etnicitet	ethnicity	0	0	1	0
etnicitet	ethnic	0	0	1	0
skogen	woods	0	0	1	0
skogen	forest	0	0	1	0
skilja	seperate	0	0	1	0
skilja	differ; differentiate	0	0	1	0
skilja	separate	0	0	1	1
höjdes	increased	0	0	1	0
höjdes	was raised	0	0	1	0
höjder	altitudes	0	0	1	0
höjder	heights	0	0	1	0
american	american	0	0	1	0
höjden	hojde	0	0	1	0
höjden	height	0	0	1	0
kung	king	0	0	1	1
skiljs	separated	0	0	1	0
skiljs	separate	0	0	1	0
utvecklats	developed	0	0	1	0
synen	the view	0	0	1	0
synen	sight	0	0	1	0
etiska	ehtical	0	0	1	0
etiska	codes	0	0	1	0
elden	fire	0	0	1	0
elden	the fire	0	0	1	0
fabriker	plants	0	0	1	0
fabriker	factories	0	0	1	0
helsingborgs	helsing borg	0	0	1	0
helsingborgs	helsingborg's	0	0	1	0
taggar	twig	0	0	1	0
taggar	thorn	0	0	1	0
taggar	spikes	0	0	1	0
taggar	tags	0	0	1	0
ödleblad	lizardtail	1	0	1	0
ödleblad	dleblad	1	0	1	0
ödleblad	houttuynia	1	1	0	0
ödleblad	lizard blade	1	0	1	0
ödleblad	houttuynia cordata	1	0	1	0
ödleblad	colour	1	0	1	0
ödleblad	odleblad	1	0	1	0
ödleblad	color	1	0	1	0
ödleblad	lizardleaf	1	0	1	0
ödleblad	lizard tail	1	1	0	0
ödleblad	Ödleblad	1	0	1	0
ödleblad	ödleblad	1	0	1	0
ödleblad	chameleon plant	1	1	0	0
synes	seems to	0	0	1	0
synes	apparently	0	0	1	0
synes	appears	0	0	1	0
miss	miss	0	0	1	1
rygg	dorsal	0	0	1	0
rygg	backs	0	0	1	0
rygg	back	0	0	1	1
deltagare	contestant	0	0	1	0
deltagare	participants	0	0	1	0
deltagare	participiant	0	0	1	0
nederbörd	rainfall	0	0	1	1
nederbörd	precipitation	0	0	1	0
personlighetsstörning	personality disorder	0	0	1	0
kanada	canada	0	0	1	1
kongresspartiet	congress party	0	0	1	0
kongresspartiet	indian national congress	0	0	1	0
målningen	milling	0	0	1	0
målningen	the painting	0	0	1	0
station	station	0	0	1	1
parlamentsvalet	parliament election	0	0	1	0
parlamentsvalet	election to parliament	0	0	1	0
parlamentsvalet	parliamentary elections	0	0	1	0
märktes	labeled	0	0	1	0
östberg	Östberg	0	0	1	0
östberg	ostberg	0	0	1	0
nigeria	nigeria	0	0	1	1
förstördes	destroyed	0	0	1	0
förstördes	rapids dared	0	0	1	0
förstördes	was destroyed	0	0	1	0
brittiska	british	0	0	1	0
luminositet	luminosity	0	0	1	1
brittiske	british	0	0	1	0
förebyggande	preventing	0	0	1	1
förebyggande	preventive	0	0	1	1
förebyggande	prevention	0	0	1	1
representera	represents	0	0	1	0
representera	represent	0	0	1	1
öppna	open	0	0	1	1
brittiskt	brittish	0	0	1	0
brittiskt	british	0	0	1	0
tvungen	forced	0	0	1	1
tvungen	had	0	0	1	0
tvungen	forced (to)	0	0	1	0
bildande	forming	0	0	1	0
bildande	founding	0	0	1	0
bildande	formation	0	0	1	1
brasiliens	brazil's	0	0	1	0
läggs	is	0	0	1	0
läggs	put before; submitted; put	0	0	1	0
läggs	lay	0	0	1	0
aristokratin	the aristocraty	0	0	1	0
aristokratin	aristocracy	0	0	1	0
andersson	andersson	0	0	1	0
sämsta	worst	0	0	1	0
haddock	haddock	0	0	1	0
lägga	put	0	0	1	1
lägga	add	0	0	1	0
lägga	lay	0	0	1	1
stiftelsen	foundation	0	0	1	0
linnés	linnaeus	0	0	1	0
gren	crotch	0	0	1	1
gren	branch	0	0	1	1
sekunder	seconds	0	0	1	0
sekunder	second	0	0	1	0
charlotte	charlotte	0	0	1	0
missförstånd	misunderstanding	0	0	1	1
missförstånd	misunderstandings	0	0	1	0
teslas	teslas	0	0	1	0
teslas	tesla's	0	0	1	0
genomgripande	radical	0	0	1	0
genomgripande	good	0	0	1	0
genomgripande	comprehensive; radical	0	0	1	0
medeltemperaturen	median temperature	0	0	1	0
medeltemperaturen	the average temperature	0	0	1	0
nominerad	nominate	0	0	1	0
nominerad	nominated	0	0	1	0
karl	karl	0	0	1	0
godkände	approved	0	0	1	0
genomföra	perform	0	0	1	0
genomföra	out	0	0	1	0
liberalismen	the liberalism	0	0	1	0
liberalismen	liberalism	0	0	1	0
henne	she	0	0	1	0
henne	her	0	0	1	1
liv	life	0	0	1	1
herre	lord	0	0	1	1
herre	master; lord	0	0	1	0
avseenden	respects	0	0	1	0
avseenden	regard	0	0	1	0
genomförs	conducted	0	0	1	0
genomförs	implemented	0	0	1	0
genomförs	is carried out	0	0	1	0
genomförs	carried through	0	0	1	0
genomfört	carried out	0	0	1	0
genomfört	implemented	0	0	1	0
genomfört	carried through	0	0	1	0
mexiko	mexico	0	0	1	0
logotyp	logo	0	0	1	1
logotyp	logotype	0	0	1	1
sektor	sector	0	0	1	1
kan	can be	0	0	1	0
freddie	freddie	0	0	1	0
kap	chapter	0	0	1	0
kap	cape	0	0	1	1
folkmängden	population	0	0	1	0
ledaren	leader	0	0	1	0
ledaren	conductor	0	0	1	0
användning	use	0	0	1	1
användning	use; usage	0	0	1	0
himlakroppar	celestial bodies	0	0	1	0
stå	stand	0	0	1	1
fötter	feet	0	0	1	0
fötter	on its feet	0	0	1	0
djurgårdens	djurgården's	0	0	1	0
polacker	polish	0	0	1	0
polacker	poles	0	0	1	0
företagets	the company's	0	0	1	0
företagets	the corporation's	0	0	1	0
försäljningen	gush sales	0	0	1	0
försäljningen	sales	0	0	1	0
recensioner	reviews	0	0	1	0
ingenting	nothing	0	0	1	1
jupiters	jupiter's	0	0	1	0
jupiters	jupiter	0	0	1	0
förbjudna	forbidden	0	0	1	0
förbjudna	prohibited	0	0	1	0
counterstrike	counterstrike	0	0	1	0
loggbok	log book	1	0	1	0
loggbok	journal	1	1	0	1
loggbok	analogue	1	0	1	0
loggbok	logbook	1	1	0	0
loggbok	log	1	0	1	1
muslimsk	muslim	0	0	1	1
muslimsk	muslim; muslem	0	0	1	0
svenskans	the swedish language	0	0	1	0
svenskans	swedish language	0	0	1	0
justice	justice	0	0	1	0
dröm	dream	0	0	1	1
dröm	syndrome	0	0	1	0
mullusfiskar	mullusfiskar (fish)	1	0	1	0
mullusfiskar	mullets	1	0	1	0
mullusfiskar	don't know what it is except for a kind of fish	1	0	1	0
mullusfiskar	fish	1	0	1	0
mullusfiskar	goatfish	1	1	0	0
mullusfiskar	mullusfiskar	1	0	1	0
mullusfiskar	red mullet	1	0	1	0
mullusfiskar	admit	1	0	1	0
mullusfiskar	mullisfiskar (fish)	1	0	1	0
mullusfiskar	accept	1	0	1	0
mullusfiskar	allow	1	0	1	0
mullusfiskar	perch fish	1	1	0	0
mullusfiskar	mullet	1	0	1	0
mullusfiskar	goatfishes	1	0	1	0
humanistiska	humane	0	0	1	0
humanistiska	humanistic	0	0	1	0
humanistiska	humanist	0	0	1	0
ikon	icon	0	0	1	1
darwin	darwin	0	0	1	0
blått	blue	0	0	1	0
somalia	somalia	0	0	1	0
grön	green	0	0	1	1
utrikes	foreign	0	0	1	1
måne	moon	0	0	1	1
återkommande	recurring	0	0	1	1
upphovsrätten	copyright	0	0	1	0
alexander	alexander	0	0	1	0
östfronten	eastern front	0	0	1	0
östfronten	the east front	0	0	1	0
östfronten	eastern	0	0	1	0
avsaknaden	absence	0	0	1	0
baháí	baha'i	0	0	1	0
baháí	bahá'í	0	0	1	0
vilken	what	0	0	1	1
vilken	which	0	0	1	1
vilket	which	0	0	1	1
lägsta	lowest	0	0	1	0
lägsta	minimum	0	0	1	0
x	x	0	0	1	0
tolkiens	tolkien's	0	0	1	0
tolkiens	tolkien	0	0	1	0
grunden	base	0	0	1	0
grunden	basis	0	0	1	0
spaniens	spain's	0	0	1	0
stärka	enhance	0	0	1	0
stärka	strong	0	0	1	0
stärka	strengthen; bolster	0	0	1	0
bakgrund	background	0	0	1	1
bakgrund	bakground	0	0	1	0
tidigare	earlier	0	0	1	0
tidigare	before	0	0	1	0
kanarieöarna	canary islands	0	0	1	0
kanarieöarna	the canary islands	0	0	1	0
grunder	bases	0	0	1	0
flyter	float	0	0	1	0
flyter	flows	0	0	1	0
chefen	head	0	0	1	0
chefen	commendant; commander	0	0	1	0
åsikten	the opinion	0	0	1	0
åsikten	view	0	0	1	0
pictures	pictures	0	0	1	0
påstås	claimed	0	0	1	0
påstås	(been) said	0	0	1	0
påstås	allegedly	0	0	1	0
påstår	states	0	0	1	0
påstår	claims	0	0	1	0
påstår	asserts	0	0	1	0
filmen	the movie	0	0	1	0
filmen	film	0	0	1	0
åsikter	opinions	0	0	1	0
produkten	product	0	0	1	0
produkten	the result	0	0	1	0
sålts	sold	0	0	1	0
förbli	remain	0	0	1	1
chansen	chances	0	0	1	0
chansen	chance	0	0	1	0
allvar	earnest	0	0	1	0
allvar	serious	0	0	1	0
likhet	resemblance	0	0	1	1
likhet	similar	0	0	1	0
likhet	like	0	0	1	0
gudomlig	divine	0	0	1	1
atmosfären	atmosphere	0	0	1	0
atmosfären	the atmosphere	0	0	1	0
genre	genre	0	0	1	1
produkter	products	0	0	1	0
league	league	0	0	1	0
lejonet	havskattfskar	0	0	1	0
lejonet	the lion	0	0	1	0
lejonet	lion	0	0	1	0
anor	ancestry	0	0	1	1
anor	lineage; ancestry	0	0	1	0
boende	resident	0	0	1	1
boende	housing	0	0	1	0
boende	accommodation	0	0	1	0
viljan	will	0	0	1	0
viljan	te will	0	0	1	0
slavar	slaves	0	0	1	0
kyrkliga	religious	0	0	1	0
kyrkliga	from the church	0	0	1	0
kyrkliga	church	0	0	1	0
bott	lived	0	0	1	0
bott	lived in	0	0	1	0
städerna	city ​​limits	0	0	1	0
städerna	urban	0	0	1	0
städerna	the towns	0	0	1	0
evolutionsteorin	theory of evolution	0	0	1	0
sägs	said (to be)	0	0	1	0
sägs	said	0	0	1	0
betydde	meant	0	0	1	0
betydde	ment	0	0	1	0
scientologikyrkan	the church of scientology	0	0	1	0
scientologikyrkan	church of scientology	0	0	1	0
säga	say	0	0	1	1
linux	linux	0	0	1	0
sokrates	socrates	0	0	1	1
sokrates	sokrates	0	0	1	0
planeter	planets	0	0	1	0
skydd	protection	0	0	1	1
merparten	most	0	0	1	0
merparten	the majority	0	0	1	0
merparten	larger part	0	0	1	0
arsenal	arsenal	0	0	1	1
minskade	minimum period	0	0	1	0
minskade	was reduced	0	0	1	0
minskade	decreased	0	0	1	0
söker	searches	0	0	1	0
söker	seek	0	0	1	0
söker	seeks out	0	0	1	0
enheten	the unit	0	0	1	0
enheten	unit	0	0	1	0
enheter	units	0	0	1	0
kuster	coasts	0	0	1	0
konsensus	consensus	0	0	1	0
gestalt	character	0	0	1	1
gestalt	figure	0	0	1	1
walter	walter	0	0	1	0
fåglarna	the birds	0	0	1	0
fåglarna	birds	0	0	1	0
återfinns	found	0	0	1	0
återfinns	is rediscovered	0	0	1	0
handlingen	hand-writing	0	0	1	0
handlingen	the plot	0	0	1	0
handlingen	the story	0	0	1	0
budgeten	budget	0	0	1	0
budgeten	the budget	0	0	1	0
anthony	anthony	0	0	1	0
livet	the life	0	0	1	0
livet	life	0	0	1	0
anspråk	claims	0	0	1	0
anspråk	claim	0	0	1	1
delades	shared	0	0	1	0
delades	divided	0	0	1	0
delades	split	0	0	1	0
socialism	socialism	0	0	1	1
match	game	0	0	1	1
match	match	0	0	1	1
hegel	hegel	0	0	1	0
diktator	dictator	0	0	1	1
diktator	siktador	0	0	1	0
guide	guide	0	0	1	1
slutar	ends	0	0	1	0
slutar	end	0	0	1	0
slutat	ended	0	0	1	0
slutat	left	0	0	1	0
kategorikvinnor	category women	0	0	1	0
nationalitet	nationality	0	0	1	1
klippiga	rocky	0	0	1	0
lagar	laws	0	0	1	0
framåt	forward	0	0	1	1
framåt	forth	0	0	1	1
kombineras	combined	0	0	1	0
staffan	staffan	0	0	1	0
kombinerat	combined	0	0	1	0
grant	word	0	0	1	0
borgerliga	bourgeois	0	0	1	0
borgerliga	conservative	0	0	1	0
deltagande	participation	0	0	1	1
sammanlagt	a total of	0	0	1	0
sammanlagt	total	0	0	1	0
sammanlagt	totaly	0	0	1	0
demokratin	the democracy	0	0	1	0
demokratin	democracy	0	0	1	0
kombinerad	combined	0	0	1	1
grand	grand	0	0	1	0
inledde	started	0	0	1	0
inledde	launched	0	0	1	0
folkslag	kind of people	0	0	1	0
folkslag	peoples	0	0	1	0
kungahuset	royal family	0	0	1	0
kungahuset	royal house	0	0	1	0
anklagats	accused	0	0	1	0
kommunicera	communicate	0	0	1	1
kommunicera	communicating	0	0	1	0
seglade	sailed	0	0	1	0
armenien	armenien	0	0	1	0
armenien	armenian	0	0	1	0
armenien	armenia	0	0	1	1
svealand	svealand	0	0	1	0
ohälsa	disorders	0	0	1	0
fatta	make	0	0	1	0
fatta	to make	0	0	1	0
kurdisk	kurdish	0	0	1	1
cruz	cruz	0	0	1	0
flygplan	aircraft	0	0	1	1
flygplan	airplane	0	0	1	1
nutid	present day	0	0	1	0
nutid	present	0	0	1	0
diagnosen	diagnosis	0	0	1	0
diagnosen	the diagnose	0	0	1	0
innersta	innermost	0	0	1	0
innersta	inner	0	0	1	0
tillverkning	production	0	0	1	1
österrikiska	austrian	0	0	1	0
hotell	hotel	0	0	1	1
njurarna	the kidneys	0	0	1	0
njurarna	kidney	0	0	1	0
tortyr	torture	0	0	1	1
skal	shell	0	0	1	1
skal	skin	0	0	1	1
fredliga	peacefull	0	0	1	0
fredliga	peaceful	0	0	1	0
romerskkatolska	roman catholic	0	0	1	0
schack	schack	1	0	1	0
schack	zircon	1	0	1	0
schack	shack	1	0	1	0
schack	chess	1	1	0	1
schack	performance	1	0	1	0
schack	execution	1	0	1	0
schack	check	1	0	1	1
uppfinnare	inventor	0	0	1	1
kallblod	cold blood	0	0	1	0
kallblod	cold blooded	0	0	1	0
kallblod	draught horse	0	0	1	0
väckt	brought	0	0	1	0
väckt	awaken	0	0	1	0
väckt	woken	0	0	1	0
taiwan	taiwan	0	0	1	0
lik	similar	0	0	1	1
lik	alike	0	0	1	0
folkomröstning	referendum	0	0	1	1
$	s	0	0	1	0
ansåg	thought	0	0	1	0
ansåg	found	0	0	1	0
ansåg	considered	0	0	1	0
nikki	nikki	0	0	1	0
håret	hair	0	0	1	0
håret	the hair	0	0	1	0
barack	barack	0	0	1	0
barack	barracks	0	0	1	1
intäkterna	the revenues	0	0	1	0
intäkterna	proceeds	0	0	1	0
intäkterna	the revenue	0	0	1	0
varuhus	warehouse	0	0	1	0
varuhus	department store	0	0	1	1
egenskap	trait	0	0	1	1
egenskap	ability	0	0	1	0
egenskap	seeks	0	0	1	0
djup	deep	0	0	1	1
marco	marco	0	0	1	0
producerats	produced	0	0	1	0
producerats	produced (by)	0	0	1	0
döpte	renamed	0	0	1	0
döpte	baptized	0	0	1	1
kulturen	culture	0	0	1	0
kulturen	the culture	0	0	1	0
avgör	determines	0	0	1	0
avgör	decides	0	0	1	0
avgör	avor	0	0	1	0
kulturer	cultures	0	0	1	0
gitarristen	the guitarist	0	0	1	0
gitarristen	guitarists	0	0	1	0
game	game	0	0	1	0
baserade	based	0	0	1	0
unga	young	0	0	1	0
immigranter	immigrants	0	0	1	0
innan	before	0	0	1	1
releasedatum	release date	0	0	1	0
dylikt	such	0	0	1	0
infektion	infection	0	0	1	1
criss	criss	0	0	1	0
gandhis	gandhi's	0	0	1	0
gandhis	gandhi	0	0	1	0
terminologi	terminology	0	0	1	1
judar	jews	0	0	1	0
asiatiska	asiatic	0	0	1	0
asiatiska	asian	0	0	1	0
donna	donna	0	0	1	0
idé	regard	0	0	1	0
idé	ide	0	0	1	0
tolkats	interpretation	0	0	1	0
tolkats	interpret	0	0	1	0
tolkats	interpreted	0	0	1	0
kommenterade	comment	0	0	1	0
kommenterade	commented	0	0	1	0
byggnader	buildings	0	0	1	0
byggnader	structures	0	0	1	0
pierre	pierre	0	0	1	0
economic	economic	0	0	1	0
economic	ecomomic	0	0	1	0
publiceringen	the publication	0	0	1	0
publiceringen	publishing	0	0	1	0
publiceringen	publication	0	0	1	0
syndrom	syndrome	0	0	1	1
syndrom	syndrom	0	0	1	0
bäste	best	0	0	1	0
bästa	the best	0	0	1	0
bästa	best	0	0	1	0
skapat	created	0	0	1	0
regissör	director	0	0	1	1
förväntas	expected	0	0	1	0
hellström	hellström	0	0	1	0
hellström	hellstrom	0	0	1	0
vilda	wild	0	0	1	0
skapar	creates	0	0	1	0
skapas	creates	0	0	1	0
bestämmer	estammer	0	0	1	0
bestämmer	determines	0	0	1	0
bestämmer	decide	0	0	1	0
faktorn	factor	0	0	1	0
uppträdde	appeared	0	0	1	0
uppträdde	perform	0	0	1	0
uppträdde	occurred	0	0	1	0
spänner	spanner	0	0	1	0
spänner	span	0	0	1	0
slash	slash	0	0	1	0
föreslog	suggested	0	0	1	0
föreslog	propose	0	0	1	0
enormt	gigantic	0	0	1	0
enormt	fusionenormously	0	0	1	0
enormt	enormously	0	0	1	0
sarajevo	sarajevo	0	0	1	0
run	run	0	0	1	0
steg	rose	0	0	1	0
steg	step	0	0	1	1
rum	(took) place	0	0	1	0
rum	room	0	0	1	1
depolarisering		1	0	1	0
depolarisering	de-polarizing	1	0	1	0
depolarisering	nikolayevich	1	0	1	0
depolarisering	depolarisation	1	0	1	0
depolarisering	depolarization	1	1	0	0
depolarisering	nikolaevich	1	0	1	0
sten	stone	0	0	1	1
mellankrigstiden	interwar period	0	0	1	0
mellankrigstiden	time between the wars	0	0	1	0
mellankrigstiden	interwar years	0	0	1	0
fördrevs	was banished	0	0	1	0
fördrevs	ford described	0	0	1	0
fördrevs	driven away	0	0	1	0
offside	offside	0	0	1	1
benfica	benfica	0	0	1	0
järnvägen	railroad	0	0	1	0
järnvägen	rail	0	0	1	0
myndighet	authoroty	0	0	1	0
myndighet	authority	0	0	1	1
linjen	the line	0	0	1	0
linjen	line	0	0	1	0
etablerade	established	0	0	1	0
överlevde	survived	0	0	1	0
fysiologiska	physiological	0	0	1	0
refererar	refer (to)	0	0	1	0
refererar	references	0	0	1	0
refererar	reference	0	0	1	0
skånes	scania's	0	0	1	0
skånes	scania	0	0	1	0
linjer	routes	0	0	1	0
linjer	lines	0	0	1	0
edvard	edvard	0	0	1	0
edvard	edward	0	0	1	0
sjögren	sjögren	0	0	1	0
block	block	0	0	1	1
ida	ida	0	0	1	0
samlas	together	0	0	1	0
reaktorer	reactors	0	0	1	0
revolutionär	revolutionary	0	0	1	1
revolutionär	revolutions	0	0	1	0
närvaro	attendance	0	0	1	1
närvaro	presence	0	0	1	1
västmakterna	western powers	0	0	1	0
befolkningens	population	0	0	1	0
befolkningens	population's	0	0	1	0
sprida	spread	0	0	1	1
fokuserade	concentrated	0	0	1	0
fokuserade	focused	0	0	1	0
framfördes	were	0	0	1	0
framfördes	framfordes	0	0	1	0
ligga	lies	0	0	1	0
ligga	be	0	0	1	0
ligga	lie	0	0	1	1
visar	is	0	0	1	0
visar	shows	0	0	1	1
visas	is showed	0	0	1	0
visas	shown	0	0	1	0
visat	found	0	0	1	0
visat	shown	0	0	1	0
heritage	heritage	0	0	1	0
spridd	wide spread	0	0	1	0
spridd	widespread	0	0	1	0
spridd	spread	0	0	1	0
jonsson	jonsson	0	0	1	0
ledamot	member	0	0	1	1
ledamot	representative	0	0	1	0
strukturen	the structure	0	0	1	0
strukturen	structure	0	0	1	0
förbindelse	connections	0	0	1	0
förbindelse	connection	0	0	1	1
spektrumet	spectrum	0	0	1	0
larry	larry	0	0	1	0
strukturer	structures	0	0	1	0
strukturer	structure	0	0	1	0
bjöd	offered	0	0	1	0
bjöd	invited	0	0	1	0
drabbats	affected	0	0	1	0
drabbats	afflicted	0	0	1	0
skull	sake	0	0	1	1
ute	absent	0	0	1	0
ute	out	0	0	1	1
uppmärksammat	attention	0	0	1	0
uppmärksammat	noticed	0	0	1	0
nyval	re-election	0	0	1	0
nyval	new election	0	0	1	1
nyval	election	0	0	1	0
skuld	liability	0	0	1	0
skuld	debt	0	0	1	1
skuld	guilt	0	0	1	1
malin	maleic	0	0	1	0
malin	malin	0	0	1	0
område	area	0	0	1	1
trafikerade	traffic	0	0	1	0
trafikerade	frequent	0	0	1	0
trafikerade	trafficked	0	0	1	0
jönssonligan	jönssonligan	0	0	1	0
jönssonligan	jonssonligan	0	0	1	0
politik	politics	0	0	1	1
politik	policies	0	0	1	0
chelsea	chelsea	0	0	1	0
ligacupen	league cup	0	0	1	0
monarki	monarchy	0	0	1	1
månarna	moons	0	0	1	0
metall	metal	0	0	1	1
voltaires	voltaire	0	0	1	0
uppfyller	fulfills	0	0	1	0
igenom	through	0	0	1	1
krigets	the war's	0	0	1	0
krigets	war	0	0	1	0
sjunde	seventh	0	0	1	1
sökte	searched	0	0	1	0
musikens	music	0	0	1	0
musikens	the music's	0	0	1	0
kategori	category	0	0	1	1
klubbarna	clubs	0	0	1	0
klubbarna	the clubs	0	0	1	0
korn	korn	0	0	1	0
korn	barley	0	0	1	1
korn	grains	0	0	1	0
världsarvslista	world heritage list	0	0	1	0
rester	residue	0	0	1	0
rester	remains	0	0	1	1
rester	residues	0	0	1	0
dras	references)	0	0	1	0
dras	draw	0	0	1	0
dras	preferred	0	0	1	0
dras	make (assumptions	0	0	1	0
början	top	0	0	1	0
början	beginning	0	0	1	1
sköts	postponed; run	0	0	1	0
sköts	shot	0	0	1	0
sköts	handled	0	0	1	0
uppmärksammad	attention	0	0	1	0
uppmärksammad	come to attention	0	0	1	0
uppmärksammad	noted	0	0	1	0
uppmärksammad	noticed	0	0	1	0
william	william	0	0	1	0
drag	trait; characteristic; feature	0	0	1	0
drag	move	0	0	1	1
drag	characteristic	0	0	1	0
nödvändig	necessary	0	0	1	1
nödvändig	essential	0	0	1	0
kort	short	0	0	1	1
månens	the moon's	0	0	1	0
månens	the moons	0	0	1	0
månens	moon	0	0	1	0
jagar	hunts	0	0	1	0
jagar	hunting	0	0	1	0
börjar	starts	0	0	1	0
börjar	start	0	0	1	0
börjar	starts to	0	0	1	0
börjat	started	0	0	1	0
börjat	begun to	0	0	1	0
börjat	begun	0	0	1	1
kors	cross	0	0	1	1
samarbetade	collaborated	0	0	1	0
samarbetade	collaboration	0	0	1	0
värmland	wermlandia	0	0	1	0
värmland	varmland	0	0	1	0
värmland	värmland	0	0	1	0
förbudet	ban	0	0	1	0
förbudet	the union	0	0	1	0
dvd	dvd	0	0	1	0
årliga	annual	0	0	1	0
tunga	heavy	0	0	1	0
tunga	tongue	0	0	1	1
heath	heath	0	0	1	0
åriga	-year	0	0	1	0
åriga	year	0	0	1	0
säsong	season	0	0	1	1
folkliga	popular	0	0	1	0
folkliga	folk	0	0	1	0
tungt	heavy	0	0	1	1
svt	svt	0	0	1	0
vägnätet	road network	0	0	1	0
skyskrapor	high rise buildings; sky scrapers	0	0	1	0
skyskrapor	skyscrapers	0	0	1	0
stones	stones	0	0	1	0
stones	sone	0	0	1	0
bonniers	bonnier's	0	0	1	0
bonniers	bonniers	0	0	1	0
placera	position	0	0	1	1
placera	place	0	0	1	1
frigörs	released	0	0	1	0
frigörs	is released	0	0	1	0
katt	cat	0	0	1	1
ge	to give	0	0	1	0
ge	give	0	0	1	1
ga	ga	0	0	1	0
go	go	0	0	1	0
gm	by	0	0	1	0
kate	kate	0	0	1	0
baron	baron	0	0	1	1
möttes	met	0	0	1	0
toppar	(that) peaks	0	0	1	0
toppar	tops	0	0	1	0
toppar	peak	0	0	1	0
kräver	requires	0	0	1	0
skildras	is depicted	0	0	1	0
skildras	depicted	0	0	1	0
wave	wave	0	0	1	0
gärna	i'd love to	0	0	1	0
gärna	readily	0	0	1	1
rinner	running	0	0	1	0
rinner	flow	0	0	1	0
rinner	flows	0	0	1	0
kommunismen	communism	0	0	1	0
vätska	fluid	0	0	1	1
vätska	liquid	0	0	1	1
folkräkningen	census	0	0	1	0
folkräkningen	the census	0	0	1	0
michael	michael	0	0	1	0
ryan	ryan	0	0	1	0
världskriget	world war	0	0	1	0
utbredning	distribution	0	0	1	1
utbredning	distrubution	0	0	1	0
tidszoner	time zones	0	0	1	0
stift	pin	0	0	1	1
stift	diocese	0	0	1	1
akut	acute	0	0	1	1
akut	urgent	0	0	1	0
lämna	leave	0	0	1	1
lämna	supply	0	0	1	0
socialdemokratiska	socialists	0	0	1	0
socialdemokratiska	social democratic	0	0	1	0
ordspråk	saying	0	0	1	0
ordspråk	proverbs	0	0	1	0
ordspråk	proverb	0	0	1	1
zh	zh	0	0	1	0
derivator	derivative	0	0	1	0
derivator	derivatives	0	0	1	0
mussolinis	mussolini's	0	0	1	0
mussolinis	mussolini	0	0	1	0
honan	the female	0	0	1	0
honan	female	0	0	1	0
geologiska	geological	0	0	1	0
visserligen	certainly	0	0	1	1
visserligen	although	0	0	1	0
direkta	direct	0	0	1	0
intervjuer	interviews	0	0	1	0
gå	go	0	0	1	1
singapores	singapores	0	0	1	0
singapores	singapore's	0	0	1	0
geologiskt	geologically	0	0	1	0
geologiskt	geological	0	0	1	0
idéer	ideas	0	0	1	0
kinas	china's	0	0	1	0
kinas	kinase	0	0	1	0
kinas	chinas	0	0	1	0
kröntes	been crowned	0	0	1	0
kröntes	crowned	0	0	1	0
hansson	hansson	0	0	1	0
polen	poland	0	0	1	1
polen	pole	0	0	1	0
företräder	preferred trades	0	0	1	0
företräder	representing	0	0	1	0
genombrott	breakthrough	0	0	1	1
cell	cell	0	0	1	1
experiment	experiment	0	0	1	1
avancerade	advanced	0	0	1	0
valen	the elections	0	0	1	0
valen	elections	0	0	1	0
gamla	ancient	0	0	1	0
gamla	old	0	0	1	0
utrikespolitiken	foreign policy	0	0	1	0
utrikespolitiken	the foreign policy	0	0	1	0
invigdes	inaugurated	0	0	1	0
bindande	binding	0	0	1	1
innerstaden	inner city	0	0	1	0
orsaker	causes	0	0	1	0
eminem	eminem	0	0	1	0
vreeswijk	vreeswijk	0	0	1	0
vreeswijk	cohen	0	0	1	0
uppgick	total	0	0	1	0
uppgick	was	0	0	1	0
ökenråttor	known	1	0	1	0
ökenråttor	gerbil	1	1	0	0
ökenråttor	ökenrättor	1	0	1	0
ökenråttor	Ökenråttor	1	0	1	0
ökenråttor	famous	1	0	1	0
ökenråttor	gherbils	1	1	0	0
ökenråttor	desert rats	1	1	0	0
ökenråttor	Ökenrättor	1	0	1	0
ökenråttor	gerbils; desert rats	1	0	1	0
ökenråttor	gerbils	1	1	0	0
ökenråttor	okenrattor	1	1	0	0
ryska	russian	0	0	1	1
orsaken	reason	0	0	1	0
orsaken	cause	0	0	1	0
innebandy	floorball	0	0	1	0
integritet	integrity	0	0	1	1
känslor	music	0	0	1	0
känslor	feelings	0	0	1	0
utövar	exercises	0	0	1	0
utövar	carrying	0	0	1	0
utövar	exercise	0	0	1	0
biologi	biology	0	0	1	1
chans	chances	0	0	1	0
chans	chance	0	0	1	1
chans	chanse	0	0	1	0
utövas	is practised	0	0	1	0
utövas	exerted	0	0	1	0
utövas	exercised	0	0	1	0
ateism	atheism	0	0	1	1
ingå	be a part	0	0	1	0
ingå	include	0	0	1	0
ingå	be included in	0	0	1	0
dopamin	dopamine	0	0	1	0
uppfinningar	inventions	0	0	1	0
crazy	crazy	0	0	1	0
innebörden	meaning	0	0	1	0
innebörden	the significance	0	0	1	0
avsedda	aimed	0	0	1	0
avsedda	for	0	0	1	0
avsedda	intended	0	0	1	0
berättade	told	0	0	1	1
våldsam	violent	0	0	1	1
vuxen	adult	0	0	1	1
italienska	italian	0	0	1	1
berättelserna	the stories	0	0	1	0
berättelserna	stories	0	0	1	0
berättelserna	tales; stories	0	0	1	0
genetiska	genetic	0	0	1	0
français	francais	0	0	1	0
français	public	0	0	1	0
personen	person	0	0	1	0
personen	the person	0	0	1	0
genetiskt	genetically	0	0	1	0
genetiskt	genetic	0	0	1	0
coldplay	coldplay	0	0	1	0
kunde	could	0	0	1	1
personer	person	0	0	1	0
personer	people	0	0	1	1
personer	persons	0	0	1	0
oktober	october	0	0	1	1
intäkter	revenues	0	0	1	0
intäkter	incomes	0	0	1	0
råd	advice	0	0	1	1
råd	council	0	0	1	1
sjunger	sings	0	0	1	0
sjunger	singing	0	0	1	0
starten	the start	0	0	1	0
starten	start	0	0	1	0
präglats	been characterized	0	0	1	0
präglats	been marked	0	0	1	0
präglats	marked	0	0	1	0
about	about	0	0	1	0
uppstår	occur	0	0	1	0
balkanhalvön	balkans	0	0	1	0
balkanhalvön	balkan peninsula	0	0	1	0
lagförslag	bill	0	0	1	1
lagförslag	lagforslag	0	0	1	0
invigningen	inauguration	0	0	1	0
invigningen	the opening	0	0	1	0
huxley	huxley	0	0	1	0
överbefälhavare	commander-in-chief	0	0	1	1
överbefälhavare	overbefalhaare	0	0	1	0
överbefälhavare	supreme commander	0	0	1	0
misslyckades	failed	0	0	1	0
turkiets	turkey's	0	0	1	0
turkiets	turkeys	0	0	1	0
debutalbum	debut album	0	0	1	0
präst	priest	0	0	1	1
godkännas	approved	0	0	1	0
godkännas	pass on	0	0	1	0
godkännas	be approved	0	0	1	0
mottagaren	the receiver	0	0	1	0
mottagaren	the recipient	0	0	1	0
mottagaren	receiver	0	0	1	0
tillåter	allows	0	0	1	0
tillåter	allow	0	0	1	0
tillåtet	distillate	0	0	1	0
tillåtet	allowed	0	0	1	0
spåras	stored	0	0	1	0
spåras	trace	0	0	1	0
kenny	kenny	0	0	1	0
liknade	similar	0	0	1	0
liknade	looked like	0	0	1	0
halloween	halloween	0	0	1	0
jämföra	compare	0	0	1	1
dominans	dominant	0	0	1	0
dominans	dominance	0	0	1	1
geomorfologi	geomorphology	1	1	0	1
geomorfologi	stability	1	0	1	0
geomorfologi	stable	1	0	1	0
jämfört	compared to last	0	0	1	0
jämfört	compared	0	0	1	0
jämfört	compared (to)	0	0	1	0
studioalbum	studio album	0	0	1	0
läsning	read	0	0	1	1
läsning	reading	0	0	1	1
förstod	understood	0	0	1	0
talat	spoken	0	0	1	0
talat	spoke	0	0	1	0
talas	spoken	0	0	1	0
talas	is spoken	0	0	1	0
talar	speaks	0	0	1	0
talar	talk	0	0	1	0
talar	speak	0	0	1	0
romantikens	the romanticism	0	0	1	0
romantikens	romanticism	0	0	1	0
romantikens	romantick	0	0	1	0
bönder	farmers	0	0	1	0
georg	georgian	0	0	1	0
georg	georg	0	0	1	0
löften	promises	0	0	1	0
översättas	translated	0	0	1	0
översättas	be translated	0	0	1	0
översättas	translated (to)	0	0	1	0
sovjetunionen	the soviet union	0	0	1	0
sovjetunionen	soviet union	0	0	1	0
ferdinand	ferdinand	0	0	1	0
kronprinsen	crown prince	0	0	1	0
kronprinsen	the crown prince	0	0	1	0
oroligheter	unrest	0	0	1	0
fara	danger	0	0	1	1
uttalet	the pronounciation	0	0	1	0
uttalet	pronunciation	0	0	1	0
ronald	ronald	0	0	1	0
fart	speed	0	0	1	1
fart	off	0	0	1	0
fars	father's	0	0	1	0
fars	father	0	0	1	0
ringde	called	0	0	1	0
västberlin	west berlin	0	0	1	0
beskrivningen	description	0	0	1	0
reagerar	react	0	0	1	0
reagerar	reacts	0	0	1	0
möjligheter	mojligheter	0	0	1	0
möjligheter	potential	0	0	1	0
övriga	other	0	0	1	0
övriga	others	0	0	1	0
solsystemets	solar system	0	0	1	0
möjligheten	the ability	0	0	1	0
möjligheten	possibility	0	0	1	0
möjligheten	the possibility	0	0	1	0
väte	hydrogen	0	0	1	1
encyclopedia	encyclopedia	0	0	1	0
kungliga	royal	0	0	1	0
innebär	means	0	0	1	0
innebär	mean	0	0	1	0
socken	parish	0	0	1	1
obelix	obelix	0	0	1	0
timmar	hours	0	0	1	0
presidenter	presidents	0	0	1	0
presidenter	president	0	0	1	0
offentliga	public	0	0	1	0
månad	month	0	0	1	1
bosättningar	settlements	0	0	1	0
bosättningar	bosattningar	0	0	1	0
presidenten	president	0	0	1	0
presidenten	the president	0	0	1	0
månar	moons	0	0	1	0
närhet	close	0	0	1	0
närhet	proximity	0	0	1	0
närhet	closeness	0	0	1	1
verklighet	true	0	0	1	0
verklighet	reality	0	0	1	1
belopp	amounts	0	0	1	0
belopp	amount	0	0	1	1
belopp	sum	0	0	1	1
begick	commited	0	0	1	0
begick	committed	0	0	1	0
kyrkor	churche	0	0	1	0
kyrkor	churches	0	0	1	0
insekter	insects	0	0	1	0
tätbefolkade	densely populated	0	0	1	0
tätbefolkade	populated	0	0	1	0
allting	everything	0	0	1	1
filosofiska	philosophical	0	0	1	0
naturgas	natural gas	0	0	1	1
konserten	the concert	0	0	1	0
konserten	concert	0	0	1	0
zagreb	capital of croatia	0	0	1	0
zagreb	zagreb	0	0	1	0
säljer	sells	0	0	1	0
lån	loan	0	0	1	1
restauranger	restaurants	0	0	1	0
restauranger	restaurant	0	0	1	0
låt	let	0	0	1	0
låt	methacrylate	0	0	1	0
låt	song	0	0	1	1
fördel	advantageously	0	0	1	0
fördel	advantage	0	0	1	1
front	front	0	0	1	1
konserter	conserts	0	0	1	0
konserter	concerts	0	0	1	0
dikt	poem	0	0	1	1
miniatyr|px|den	miniature	0	0	1	0
hunden	the dog	0	0	1	0
hunden	dog	0	0	1	0
university	university	0	0	1	0
finnas	found	0	0	1	0
finnas	exists	0	0	1	0
finnas	(be) found	0	0	1	0
nordirland	north ireland	0	0	1	0
nordirland	northern	0	0	1	0
stöd	support	0	0	1	1
mode	fashion	0	0	1	1
mode	mode	0	0	1	1
förändring	alteration	0	0	1	1
förändring	change	0	0	1	1
modo	modo	0	0	1	0
stadsparken	city park	0	0	1	0
stadsparken	stadsparken	0	0	1	0
stadsparken	city ​​park	0	0	1	0
skog	wood	0	0	1	1
skog	forest	0	0	1	1
globe	globe	0	0	1	0
åtskilda	separated	0	0	1	0
åtskilda	segregated	0	0	1	0
åtskilda	separate	0	0	1	0
stiger	rises	0	0	1	0
stiger	rising	0	0	1	0
osmanerna	ottoman turks	0	0	1	0
osmanerna	ottomans	0	0	1	0
osmanerna	osmanerna	0	0	1	0
skov	forestry	0	0	1	0
skov	episode	0	0	1	0
skov	relapse	0	0	1	0
skor	shoe	0	0	1	0
skor	shoes	0	0	1	1
special	special	0	0	1	0
flyr	flees	0	0	1	0
flyr	escapes	0	0	1	0
kärnkraftverk	nuclear power plant	0	0	1	0
kärnkraftverk	nuclear powerplant	0	0	1	0
entertainment	entertainment	0	0	1	0
huvudstad	capital city	0	0	1	0
huvudstad	capital	0	0	1	1
samarbetar	cooperates	0	0	1	0
samarbetar	collaborates	0	0	1	0
samarbetar	cooperate	0	0	1	0
samarbetat	collaborated	0	0	1	0
samarbetat	collobrated	0	0	1	0
max	max	0	0	1	0
solsystem	solar system	0	0	1	1
utgör	constitutes	0	0	1	0
utgör	make up	0	0	1	0
sällskapet	society	0	0	1	0
sällskapet	the company	0	0	1	0
vinter	winter	0	0	1	1
omfatta	cover	0	0	1	1
torres	torres	0	0	1	0
kropp	body	0	0	1	1
bilder	images	0	0	1	0
bilder	pictures	0	0	1	1
lycka	happiness	0	0	1	1
lycka	good luck	0	0	1	0
lida	sheath	0	0	1	0
lida	suffer	0	0	1	1
fastställdes	confirmed	0	0	1	0
fastställdes	set	0	0	1	0
fastställdes	laid down that	0	0	1	0
bilden	image	0	0	1	0
bilden	the image	0	0	1	0
döda	dead	0	0	1	0
kommunala	local	0	0	1	0
kommunala	municipal	0	0	1	0
användbar	useful	0	0	1	1
livsmedel	food	0	0	1	1
banor	paths	0	0	1	0
banor	line	0	0	1	0
times	times	0	0	1	0
strida	conflict	0	0	1	1
strida	fight	0	0	1	1
tigrar	tigers	0	0	1	0
austin	austin	0	0	1	0
tvungna	forced	0	0	1	0
tvungna	forced to	0	0	1	0
praxis	practice	0	0	1	0
riksdagsvalet	parliamentary election	0	0	1	0
riksdagsvalet	election to parliament	0	0	1	0
riksdagsvalet	parliamentary elections	0	0	1	0
evans	mr. evans	0	0	1	0
evans	evans	0	0	1	0
förenade	united	0	0	1	0
möts	meet	0	0	1	0
möts	meets	0	0	1	0
mött	faced	0	0	1	0
mött	met	0	0	1	0
kategorihedersdoktorer	category of honorary degrees	0	0	1	0
förekomma	occur	0	0	1	1
förekomma	be found	0	0	1	1
maurice	maurice	0	0	1	0
attack	attack	0	0	1	1
boken	paper	0	0	1	0
boken	the book	0	0	1	0
dygnet	day	0	0	1	0
infaller	no cells	0	0	1	0
infaller	falls	0	0	1	0
final	finite	0	0	1	0
final	final	0	0	1	1
rumänska	romanian	0	0	1	1
viktor	viktor	0	0	1	0
belgiska	belgian	0	0	1	0
hasch	hashish	0	0	1	1
emellertid	however	0	0	1	1
höftledsgrop	hoftledsgrop	1	0	1	0
höftledsgrop	concave joint surface	1	0	1	0
höftledsgrop	mineral	1	0	1	0
höftledsgrop	acetabulum	1	1	0	0
höftledsgrop	hip pit	1	0	1	0
höftledsgrop	hip bone	1	1	0	0
höftledsgrop	hip joint	1	0	1	0
höftledsgrop	aetabulum	1	0	1	0
höftledsgrop	hip joint fossa	1	0	1	0
höftledsgrop	minerals	1	0	1	0
höftledsgrop	ores	1	0	1	0
styrelseskick	form of government	0	0	1	0
styrelseskick	government	0	0	1	0
lista	list	0	0	1	1
hushåll	household	0	0	1	1
representerade	represented	0	0	1	0
representerade	represent	0	0	1	0
ben	bone	0	0	1	1
definieras	defined	0	0	1	0
definieras	is defined	0	0	1	0
definieras	defines	0	0	1	0
definierar	defining	0	0	1	0
definierar	defines	0	0	1	0
arbetade	worked	0	0	1	0
israelisk	israeli	0	0	1	1
ber	ask	0	0	1	0
ber	asks	0	0	1	0
förlora	lose	0	0	1	1
nämnde	mentioned	0	0	1	0
nämnde	said	0	0	1	0
bet	bit	0	0	1	0
monografi	monography	1	1	0	0
monografi	monografia	1	1	0	0
monografi	every	1	0	1	0
monografi	thesis	1	0	1	0
monografi	each	1	0	1	0
monografi	monograph	1	1	0	1
lösningar	solutions	0	0	1	0
kvinnans	female	0	0	1	0
need	need	0	0	1	0
bordet	the table	0	0	1	0
bordet	desktop	0	0	1	0
varade	duration	0	0	1	0
varade	lasted	0	0	1	0
turnéer	tours	0	0	1	0
förbjöds	banned	0	0	1	0
förbjöds	forbidden	0	0	1	0
tredjedelar	thirds	0	0	1	0
visor	songs	0	0	1	0
attackerna	attacks	0	0	1	0
attackerna	the attacks	0	0	1	0
attackerna	attack	0	0	1	0
runorna	the runes	0	0	1	0
runorna	runes	0	0	1	0
jorge	jorge	0	0	1	0
beslöt	resolved	0	0	1	0
beslöt	decided	0	0	1	0
regn	rain	0	0	1	1
sats	statements	1	1	0	0
sats	covering	1	0	1	0
sats	clause	1	1	0	1
sats	sentence	1	1	0	1
sats	cover	1	0	1	0
sats	kit	1	1	1	0
sats	rate	1	0	1	1
sats	proposition	1	0	1	1
sats	statement	1	0	1	0
sats	theorem	1	0	1	1
sats	theorems; sets	1	0	1	0
sats	sets	1	0	1	0
sats	proof	1	0	1	0
sats	theorem; sets	1	1	0	0
montana	montana	0	0	1	0
genomslag	breakthrough	0	0	1	0
genomslag	impact	0	0	1	0
regi	direction	0	0	1	0
ministerrådet	minister counsellor	0	0	1	0
ministerrådet	ministers	0	0	1	0
inlärning	learning	0	0	1	1
tyskar	germans	0	0	1	0
kvällen	the evening	0	0	1	0
kvällen	evening	0	0	1	0
stjärnornas	stellar	0	0	1	0
stjärnornas	the star's	0	0	1	0
borgmästare	mayor	0	0	1	1
skogar	forests	0	0	1	0
platon	platon	0	0	1	0
platon	platonic	0	0	1	0
parker	parker	0	0	1	0
parker	parks	0	0	1	0
fiktiv	fictitious	0	0	1	1
fiktiv	fictive	0	0	1	0
tolkien	tolkien	0	0	1	0
fynden	finds; findings	0	0	1	0
fynden	findings	0	0	1	0
skedde	was	0	0	1	0
passa	take the opportunity	0	0	1	0
passa	fit	0	0	1	1
passa	match	0	0	1	0
parken	park	0	0	1	0
parken	the park	0	0	1	0
förbränning	combustion	0	0	1	1
förbränning	incineration	0	0	1	1
hade	had	0	0	1	0
hade	was	0	0	1	0
basen	became	0	0	1	0
basen	the base	0	0	1	0
basen	base	0	0	1	0
baser	bases	0	0	1	0
gemensam	joint	0	0	1	1
gemensam	common	0	0	1	1
varit	has been	0	0	1	0
varit	been	0	0	1	0
partnern	partner	0	0	1	0
partnern	the partner	0	0	1	0
aspekt	aspect	0	0	1	1
psykologin	the psyhology	0	0	1	0
psykologin	psychology	0	0	1	0
boris	boris	0	0	1	0
klassiska	classic	0	0	1	0
ställde	set	0	0	1	0
ställde	stood up	0	0	1	0
ställde	asked	0	0	1	0
omloppsbana	omloppsbana	0	0	1	0
omloppsbana	orbit	0	0	1	1
michigan	michigan	0	0	1	0
inflytelserika	influential	0	0	1	0
klassiskt	classical	0	0	1	0
klassiskt	classic	0	0	1	0
tämligen	rather	0	0	1	1
tämligen	fairly	0	0	1	1
tämligen	tamil again	0	0	1	0
århundradet	century	0	0	1	0
härstamning	lineage	0	0	1	1
härstamning	origin	0	0	1	0
härstamning	descent	0	0	1	1
gray	gray	0	0	1	0
evolution	evolution	0	0	1	1
processer	processes	0	0	1	0
mohammed	mohammed	0	0	1	0
fröken	miss	0	0	1	1
grav	tomb	0	0	1	1
grav	grave	0	0	1	1
långsamt	slowly	0	0	1	0
gran	spruce	0	0	1	1
influensa	flu	0	0	1	1
influensa	influenza	0	0	1	1
influensa	flue	0	0	1	1
riksföreståndare	regent	0	0	1	1
grad	grade	0	0	1	1
grad	rate	0	0	1	0
kvadratkilometer	square kilometer	0	0	1	0
kvadratkilometer	square kilometers	0	0	1	0
processen	process	0	0	1	0
processen	the process	0	0	1	0
upplösning	resolution; dissolution	0	0	1	0
upplösning	resolution	0	0	1	1
sydafrika	south africa	0	0	1	0
påtryckningar	pressure	0	0	1	0
påtryckningar	pressures	0	0	1	0
benämningen	label	0	0	1	0
benämningen	the name	0	0	1	0
benämningen	the designation	0	0	1	0
neutralt	neutral	0	0	1	0
landsting	county	0	0	1	0
landsting	county council	0	0	1	0
immunförsvar	immune	0	0	1	0
immunförsvar	immune defense	0	0	1	0
däribland	among them	0	0	1	0
däribland	including	0	0	1	0
förkortningar	abbreviations	0	0	1	0
stats	state's	0	0	1	0
stats	state	0	0	1	0
tenn	tin	0	0	1	1
antika	ancient	0	0	1	0
flicka	pocket	1	0	1	0
flicka	jewish	1	0	1	0
flicka	girl	1	1	1	1
havskattfiskar	catfish fish	1	0	1	0
havskattfiskar	catfish fishing	1	1	0	0
havskattfiskar	congress	1	0	1	0
havskattfiskar	havskattfskar	1	0	1	0
havskattfiskar	goatfish	1	1	0	0
havskattfiskar	anarhichadidae	1	1	0	0
havskattfiskar	catfishes	1	0	1	0
havskattfiskar	catfished	1	1	0	0
havskattfiskar	catfish	1	1	0	0
havskattfiskar	wolffish	1	1	0	0
havskattfiskar	seawolf	1	0	1	0
havskattfiskar	mullet	1	0	1	0
havskattfiskar	have duty fish	1	0	1	0
havskattfiskar	sea wolfs	1	1	0	0
havskattfiskar	ocean catfish	1	0	1	0
beräknades	were calculated	0	0	1	0
beräknades	estimated	0	0	1	0
beräknades	calculated	0	0	1	0
gotiska	gothic	0	0	1	1
staty	statue	0	0	1	1
state	state	0	0	1	0
diktatorn	the dictator	0	0	1	0
diktatorn	dictator	0	0	1	0
ken	ken	0	0	1	0
ken	bank	0	0	1	0
verksamhet	work	0	0	1	0
verksamhet	activity	0	0	1	1
sovjetiska	soviet	0	0	1	0
sovjetiska	sovjet	0	0	1	0
satsa	bet	0	0	1	0
merry	merry	0	0	1	0
jobba	work	0	0	1	1
verksam	active	0	0	1	1
verksam	effective	0	0	1	0
upprättas	established	0	0	1	0
upprättas	establish	0	0	1	0
problem	problem	0	0	1	1
problem	problems	0	0	1	0
hits	hits	0	0	1	0
reguljära	regular	0	0	1	0
synvinkel	angle	0	0	1	1
synvinkel	perspective	0	0	1	0
vulkaner	volcanos	0	0	1	0
vulkaner	volcanoes	0	0	1	0
nyare	newer	0	0	1	1
stödet	support	0	0	1	0
stödet	the support	0	0	1	0
varierade	varied	0	0	1	0
stratton	stratton	0	0	1	0
partiklar	particles	0	0	1	0
jersey	jersey	0	0	1	1
helsingfors	helsingfors	0	0	1	0
helsingfors	helsinki	0	0	1	0
jim	jim	0	0	1	0
opposition	opposition	0	0	1	1
ände	of	0	0	1	0
ände	end	0	0	1	1
kategoribrittiska	category: british	0	0	1	0
kategoribrittiska	category uk	0	0	1	0
knst	knst	0	0	1	0
leipzig	liepzig	0	0	1	0
leipzig	leipzig	0	0	1	0
johans	johan's	0	0	1	0
johans	johan	0	0	1	0
revolutionen	the revolution	0	0	1	0
revolutionen	revolution	0	0	1	0
johann	johann	0	0	1	0
johann	john	0	0	1	0
kings	kings	0	0	1	0
kings	king's	0	0	1	0
kings	king	0	0	1	0
sammanhang	connection	0	0	1	1
sammanhang	context	0	0	1	1
christer	chris	0	0	1	0
christer	christer	0	0	1	0
willy	willy	0	0	1	0
likör	cordial	1	1	0	1
likör	financing	1	0	1	0
likör	liquor	1	1	0	0
likör	liqeur	1	1	0	0
likör	liquer	1	1	0	0
likör	liqueur	1	1	0	1
sara	sara	0	0	1	0
fokusera	focus	0	0	1	1
poet	poet	0	0	1	1
poes	poe	0	0	1	0
poes	poe's	0	0	1	0
poes	poes	0	0	1	0
pontus	pontus	0	0	1	0
vinci	vinci	0	0	1	0
spanska	spanish	0	0	1	0
spaniel	spaniel	0	0	1	1
spanien	spain	0	0	1	1
skärgård	archipelago	0	0	1	1
skärgård	cutting garden	0	0	1	0
skärgård	archipelagos	0	0	1	0
hamburg	hamburger	0	0	1	0
hamburg	hamburg	0	0	1	0
bråk	brawl; fight	0	0	1	0
bråk	fights	0	0	1	0
bråk	fraction	0	0	1	1
erbjuda	offer	0	0	1	1
reaktionerna	the reactions	0	0	1	0
reaktionerna	reactions	0	0	1	0
utmärker	characterizes	0	0	1	0
utmärker	characterized	0	0	1	0
äter	eat	0	0	1	0
äter	eats	0	0	1	0
undersökte	investigated	0	0	1	0
undersökte	examined	0	0	1	0
utgjorde	made up	0	0	1	0
utgjorde	was	0	0	1	0
utgjorde	comprised; consisted of	0	0	1	0
känslig	susceptible	0	0	1	0
platons	platon's	0	0	1	0
platons	plato	0	0	1	0
platons	platos	0	0	1	0
reaktion	reaction	0	0	1	1
reaktion	reaction reaction	0	0	1	0
vilkas	volkas	0	0	1	0
vilkas	whose	0	0	1	1
rysslands	russia's	0	0	1	0
enkel	simple	0	0	1	1
enkel	plain	0	0	1	1
förklaringen	the explanation	0	0	1	0
förklaringen	statement	0	0	1	0
feber	fever	0	0	1	1
demo	demo	0	0	1	0
demo	removed	0	0	1	0
mysterium	mystery	0	0	1	1
hållning	position	0	0	1	0
hållning	attitude	0	0	1	1
hållning	entertainment	0	0	1	0
alfabetisk	alphabetical	0	0	1	1
revir	turf	0	0	1	0
revir	territory	0	0	1	1
änden	end	0	0	1	0
änden	spirit	0	0	1	0
territoriet	territory	0	0	1	0
reformationen	reformation tone	0	0	1	0
reformationen	reformation	0	0	1	0
reformationen	the reformation	0	0	1	0
gård	farm	0	0	1	0
gård	house	0	0	1	0
parti	party	0	0	1	1
parti	batch	0	0	1	0
instabil	unstable	0	0	1	1
östberlin	east berlin	0	0	1	0
campus	campus	0	0	1	0
varmed	whereby	0	0	1	1
begav	went	0	0	1	0
begav	traveled	0	0	1	0
begav	went (to)	0	0	1	0
anföll	attacked	0	0	1	0
griffon	griffon	0	0	1	0
dickens	dicken's	0	0	1	0
dickens	dickens	0	0	1	0
korrekta	correct	0	0	1	0
flygbolag	airline	0	0	1	1
flygbolag	carriers	0	0	1	0
anka	anka	0	0	1	0
anka	duck	0	0	1	1
nationens	the nation's	0	0	1	0
nationens	nation	0	0	1	0
rankas	ranks	0	0	1	0
rankas	rank	0	0	1	0
eklund	eklund	0	0	1	0
sorter	kinds	0	0	1	0
sorter	varieties	0	0	1	0
sorter	types	0	0	1	0
alperna	alps	0	0	1	1
alperna	the alps	0	0	1	0
lagring	storage	0	0	1	1
flickan	girl	0	0	1	0
flickan	the girl	0	0	1	0
grenar	branches	0	0	1	0
åtalades	was charged	0	0	1	0
åtalades	was prosecuted	0	0	1	0
åtalades	charged	0	0	1	0
i	of	0	0	1	1
i	in	0	0	1	1
övergången	transition	0	0	1	0
övergången	the transition	0	0	1	0
övergången	transformation	0	0	1	0
theodor	theodor	0	0	1	0
fläckar	stain	0	0	1	0
fläckar	stains and spots	0	0	1	0
agnostiker	agnostic	0	0	1	1
agnostiker	agnostics	0	0	1	0
onda	evil	0	0	1	0
relationer	relations	0	0	1	0
ångest	anxiety	0	0	1	1
ångest	anguish	0	0	1	1
sofia	sofia	0	0	1	0
omkom	perished	0	0	1	0
omkom	died; was killed	0	0	1	0
omkom	died	0	0	1	0
himmler	himmler	0	0	1	0
stjärnans	star's	0	0	1	0
stjärnans	the stars	0	0	1	0
stjärnans	the star's	0	0	1	0
twilight	twilight	0	0	1	0
vida	broad	0	0	1	0
vida	wide	0	0	1	0
jeff	jeff	0	0	1	0
reducera	reduce	0	0	1	1
natt	night	0	0	1	1
nato	nato	0	0	1	0
sweet	söt	0	0	1	0
titta	see	0	0	1	0
titta	watch	0	0	1	1
titta	look	0	0	1	1
bebyggelsen	building	0	0	1	0
bebyggelsen	human settlement	0	0	1	0
bebyggelsen	settlement	0	0	1	0
jesper	jesper	0	0	1	0
räknas	calculated	0	0	1	0
räknas	counted	0	0	1	0
räknas	are counted	0	0	1	0
katolska	catholic	0	0	1	0
utan	without	0	0	1	1
sanning	true	0	0	1	0
sanning	truth	0	0	1	1
underlätta	ease	0	0	1	1
underlätta	facilitate	0	0	1	1
vanligare	more common	0	0	1	0
historia	history	0	0	1	1
definitivt	permanent	0	0	1	0
definitivt	unavoidable	0	0	1	0
definitivt	definitely	0	0	1	1
historik	history	0	0	1	1
klassificering	classification	0	0	1	1
loss	off	0	0	1	0
loss	unstuck	0	0	1	1
lincoln	lincoln	0	0	1	0
lost	lost	0	0	1	0
norges	norway's	0	0	1	0
bakåt	backwards	0	0	1	1
bakåt	reverse	0	0	1	0
fernando	fernando	0	0	1	0
församlingar	parishs	0	0	1	0
församlingar	assemblies	0	0	1	0
martin	martin	0	0	1	0
auktoritära	authoritarian	0	0	1	0
regeringar	rings	0	0	1	0
regeringar	governments	0	0	1	0
jämförelser	comparison	0	0	1	0
lager	layer	0	0	1	1
våldsamma	violent	0	0	1	0
våldsamma	selection same	0	0	1	0
kolonierna	colonies	0	0	1	0
vardagliga	ordinary	0	0	1	0
vardagliga	everyday	0	0	1	0
särdrag	special features	0	0	1	0
särdrag	feature	0	0	1	1
särdrag	features	0	0	1	0
smärta	pain	0	0	1	1
pojkarna	boys	0	0	1	0
pojkarna	the boys	0	0	1	0
library	library	0	0	1	0
vardagligt	everyday	0	0	1	0
skorpan	crust	0	0	1	0
peter	peter	0	0	1	0
lagen	the law	0	0	1	0
lagen	law	0	0	1	0
moskva	moscow	0	0	1	1
skrifter	writings	0	0	1	0
jugoslaviska	jugoslavian	0	0	1	0
jugoslaviska	yugoslav	0	0	1	0
jugoslaviska	yugoslavian	0	0	1	0
spänningar	tensions	0	0	1	0
hyser	accomodates	0	0	1	0
hyser	has	0	0	1	0
hyser	holds	0	0	1	0
folkets	the people's	0	0	1	0
folkets	folkers	0	0	1	0
folkets	people	0	0	1	0
slott	castle	0	0	1	1
alliansen	the alliance	0	0	1	0
alliansen	alliance	0	0	1	0
fanns	was	0	0	1	0
skriften	no.	0	0	1	0
skriften	writings	0	0	1	0
broar	bridges	0	0	1	0
hinder	obstacle	0	0	1	1
hinder	barrier	0	0	1	0
kvarstår	remains	0	0	1	0
meddelade	stated	0	0	1	0
meddelade	announced	0	0	1	0
meddelade	informed; announced	0	0	1	0
samlades	collected	0	0	1	0
samlades	gathered	0	0	1	0
samlades	were united	0	0	1	0
journal	journal	0	0	1	1
journal	jurnal	0	0	1	0
journal	joumal	0	0	1	0
reza	reza	0	0	1	0
kromosomer	chromosomes	0	0	1	0
usas	usa:s	0	0	1	0
usas	u.s.	0	0	1	0
keramik	ceramic	0	0	1	0
keramik	ceramics	0	0	1	1
freedom	freedom	0	0	1	0
freedom	frihet	0	0	1	0
beslutade	beeslutade	0	0	1	0
beslutade	resolved	0	0	1	0
beslutade	decided	0	0	1	0
samlats	collected	0	0	1	0
samlats	solid	0	0	1	0
samlats	gathered; collected	0	0	1	0
polisens	police	0	0	1	0
polisens	the police's	0	0	1	0
troligen	probably	0	0	1	1
troligen	likely	0	0	1	0
mytologi	mythology	0	0	1	1
betydelsefulla	significant	0	0	1	0
glenn	glenn	0	0	1	0
nedan	below	0	0	1	1
nedan	hereinafter referred to as	0	0	1	0
underjordiska	underground	0	0	1	0
således	hence	0	0	1	0
således	thus	0	0	1	1
tendenser	tendencies	0	0	1	0
utility	utility	0	0	1	0
hammarby	hammarby	0	0	1	0
museum	museum	0	0	1	1
efterträddes	succeeded	0	0	1	0
realiteten	de facto	0	0	1	0
realiteten	reality	0	0	1	0
afrika	africa	0	0	1	1
heydrich	heydrich	0	0	1	0
cricket	cricket	0	0	1	0
north	north	0	0	1	0
instiftade	established	0	0	1	0
instiftade	instituted	0	0	1	0
instiftade	created	0	0	1	0
neutral	neutral	0	0	1	1
hn	hn	0	0	1	0
ho	ho	0	0	1	0
behov	necessary	0	0	1	0
hc	h.c.	0	0	1	0
hc	h.c	0	0	1	0
ha	be	0	0	1	0
ha	have	0	0	1	1
vågor	waves	0	0	1	1
he	he	0	0	1	0
samtida	contemporary	0	0	1	1
svarta	black	0	0	1	0
ljungström	ljungstrom	0	0	1	0
ljungström	ljungström	0	0	1	0
införa	introducing	0	0	1	0
införa	introduce	0	0	1	1
användningsområden	possible use	0	0	1	0
användningsområden	applications	0	0	1	0
solna	solna	0	0	1	0
fysik	physics	0	0	1	1
allierad	allied	0	0	1	1
allierad	ally	0	0	1	1
dator	computer	0	0	1	1
pippin	pippin pippin pippin	0	0	1	0
pippin	pippin	0	0	1	0
firas	celebrated	0	0	1	0
firas	celebrate	0	0	1	0
komiker	comic	0	0	1	0
komiker	comedian	0	0	1	1
isolerade	isolated	0	0	1	0
invandring	immigration	0	0	1	1
bitar	bit	0	0	1	0
bitar	pieces	0	0	1	0
beatrice	beatrice	0	0	1	0
föds	born	0	0	1	0
ordbok	glossary	0	0	1	0
ordbok	dictionary	0	0	1	1
ibland	sometimes	0	0	1	1
erik	erik	0	0	1	0
född	born	0	0	1	1
härstammar	derived	0	0	1	0
härstammar	stems	0	0	1	0
eric	eric	0	0	1	0
diego	diego	0	0	1	0
mötte	motte	0	0	1	0
mötte	met	0	0	1	0
moderaterna	the moderate	0	0	1	0
moderaterna	the moderates	0	0	1	0
moderaterna	moderates	0	0	1	0
beräkningar	calculations	0	0	1	0
speciell	specific	0	0	1	0
speciell	special	0	0	1	1
serveras	served	0	0	1	0
serveras	is served	0	0	1	0
vulkaniska	vulcanic	0	0	1	0
vulkaniska	volcanic	0	0	1	0
stat	state	0	0	1	1
hittade	found	0	0	1	0
liter	liters	0	0	1	0
dateras	dates	0	0	1	0
dateras	dated	0	0	1	0
musikvideor	music videos	0	0	1	0
framträdande	apperance	0	0	1	0
framträdande	appearance	0	0	1	1
greve	count	0	0	1	1
greve	earl	0	0	1	1
musikvideon	music video	0	0	1	0
kommersiell	commercial	0	0	1	1
stan	town	0	0	1	1
bly	led	0	0	1	0
bly	lead	0	0	1	1
stam	strain	0	0	1	0
stam	tribe	0	0	1	1
arméerna	armeerna	0	0	1	0
arméerna	armies	0	0	1	0
etiken	the ethic	0	0	1	0
etiken	ethics	0	0	1	0
succé	succes	0	0	1	0
succé	success	0	0	1	0
succé	succession	0	0	1	0
uppföljare	sequel	0	0	1	0
inser	recognize	0	0	1	0
inser	realizes	0	0	1	0
klass	grade; class	0	0	1	0
klass	class	0	0	1	1
dödlig	lethal	0	0	1	1
dödlig	mortal	0	0	1	1
alkohol	alcohol	0	0	1	1
simpson	simpson	0	0	1	0
konsumtion	consumption	0	0	1	1
hinner	reach it (in time)	0	0	1	0
hinner	have time to	0	0	1	0
hinner	time	0	0	1	0
suverän	terrific	0	0	1	0
suverän	supreme	0	0	1	0
suverän	sovereign	0	0	1	1
felaktig	incorrect	0	0	1	1
felaktig	false	0	0	1	0
felaktig	error	0	0	1	0
andre	other	0	0	1	0
protest	protest	0	0	1	1
andra	second	0	0	1	1
andra	other	0	0	1	1
fredrik	fredrik	0	0	1	0
buddy	buddy	0	0	1	0
upplagan	edition	0	0	1	0
swan	swan	0	0	1	0
kommersiellt	commercial	0	0	1	0
kulturell	cultural	0	0	1	1
bli	be	0	0	1	1
bli	become	0	0	1	1
kommersiella	commercial	0	0	1	0
passagerare	passengers	0	0	1	0
passagerare	passenger	0	0	1	1
kristendom	christianity	0	0	1	1
vasa	vasa	0	0	1	0
stormaktstiden	great power period	0	0	1	0
stormaktstiden	greatness	0	0	1	0
hemlandet	the home country	0	0	1	0
hemlandet	the homeland	0	0	1	0
examen	exam	0	0	1	1
examen	degree	0	0	1	1
disneys	disneys	0	0	1	0
disneys	disney's	0	0	1	0
disneys	disney	0	0	1	0
främst	foremost; primarily; chiefly	0	0	1	0
främst	all	0	0	1	0
främst	primarily	0	0	1	0
tätt	tight	0	0	1	1
tätt	tightly	0	0	1	0
blå	blue	0	0	1	1
blå	blah	0	0	1	0
sjö	naval	0	0	1	0
sjö	lake	0	0	1	1
chokladen	the chocolate	0	0	1	0
chokladen	chocolate	0	0	1	0
försvarsmakten	national defense	0	0	1	0
försvarsmakten	national defence	0	0	1	0
försvarsmakten	armed forces	0	0	1	0
täta	close	0	0	1	0
täta	tata	0	0	1	0
täta	seal	0	0	1	1
sexton	sixteen	0	0	1	1
dagens	current	0	0	1	0
dagens	todays	0	0	1	0
upp	up	0	0	1	1
förknippade	associated	0	0	1	0
rollfigurer	roll model	0	0	1	0
rollfigurer	role figure	0	0	1	0
rollfigurer	characters	0	0	1	0
force	force	0	0	1	0
berlins	berlin's	0	0	1	0
berlins	berlin	0	0	1	0
upplysningstiden	enlightenment	0	0	1	0
upplysningstiden	age of enlightenment	0	0	1	0
dennes	his	0	0	1	0
erövringar	conquests	0	0	1	0
avfall	waste	0	0	1	1
andré	andre	0	0	1	0
neo	neo	0	0	1	0
nej	no	0	0	1	1
kommissionen	commission	0	0	1	0
kommissionen	the commission	0	0	1	0
unescos	unesco	0	0	1	0
ned	down	0	0	1	1
ned	bottom	0	0	1	0
trodde	thought	0	0	1	0
uppträdande	performance	0	0	1	1
uppträdande	appearance	0	0	1	1
uppträdande	conduct	0	0	1	1
näsan	the nose	0	0	1	0
näsan	nose	0	0	1	0
uppdelningen	partitioning; sectionalization; division; split (-ting)	0	0	1	0
uppdelningen	splitting	0	0	1	0
uppdelningen	division	0	0	1	0
new	new	0	0	1	0
fördomar	bias	0	0	1	0
fördomar	prejudice	0	0	1	0
fördomar	prejudices	0	0	1	0
ner	bottom	0	0	1	0
romani	romani	0	0	1	0
romani	romany	0	0	1	1
romani	roma	0	0	1	0
med	with	0	0	1	1
bröts	was fractured	0	0	1	0
bröts	broke	0	0	1	0
men	but	0	0	1	1
ämnen	agents	0	0	1	0
ämnen	substances	0	0	1	1
drev	pursued	0	0	1	0
drev	drove	0	0	1	0
drev	led	0	0	1	0
vinden	the wind	0	0	1	0
vinden	wind	0	0	1	0
pedro	pedro	0	0	1	0
malmö	malmö	0	0	1	0
malmö	malmo	0	0	1	0
ämnet	substance	0	0	1	0
ämnet	subject	0	0	1	0
överföring	transfer	0	0	1	1
luther	luther	0	0	1	0
geografiskt	geographically	0	0	1	0
geografiskt	geographic	0	0	1	0
metionin	mentionin	1	0	1	0
metionin	created	1	0	1	0
metionin	methione	1	1	0	0
metionin	creation	1	0	1	0
metionin	founded	1	0	1	0
metionin	methionine	1	1	0	0
tjänst	tjanst	0	0	1	0
tjänst	service	0	0	1	1
nätet	net	0	0	1	0
nätet	the internet	0	0	1	0
dubbla	double	0	0	1	0
sju	seven	0	0	1	1
kolonier	colonies	0	0	1	0
geografiska	geographical	0	0	1	0
geografiska	spatial	0	0	1	0
dra	pulling	0	0	1	0
dra	pull; (with)draw	0	0	1	0
snabbast	fastest	0	0	1	0
magnusson	magnusson	0	0	1	0
grönland	greenland	0	0	1	1
reste	moved	0	0	1	0
reste	travelled	0	0	1	0
reste	stood	0	0	1	0
valutan	currency	0	0	1	0
rosenberg	rosenberg	0	0	1	0
stått	stood	0	0	1	0
individerna	subjects	0	0	1	0
individerna	the individuals	0	0	1	0
atlanten	atlantic	0	0	1	1
atlanten	the atlantic ocean	0	0	1	1
inleddes	started	0	0	1	0
inleddes	began	0	0	1	0
inleddes	initiated	0	0	1	0
soldat	soldier	0	0	1	1
kategorisommarvärdar	category summer hosts	0	0	1	0
prokaryoter	prokaryote	0	0	1	0
lennart	lennart	0	0	1	0
provisoriska	provisional	0	0	1	0
därmed	consequently	0	0	1	1
därmed	thus	0	0	1	0
därmed	therefore	0	0	1	0
oscar	oscar	0	0	1	0
ljus	light	0	0	1	1
nervsystemet	nervous system	0	0	1	0
nervsystemet	the nervous system	0	0	1	0
berlin	berlin	0	0	1	1
upplevde	experienced	0	0	1	0
upplevde	felt	0	0	1	0
wikipedias	wikipedia	0	0	1	0
wikipedias	wikipedias	0	0	1	0
ljud	sounds	0	0	1	0
ljud	noise	0	0	1	1
uttryckte	expressed	0	0	1	0
flora	flora	0	0	1	1
trots	although	0	0	1	0
trots	despite	0	0	1	1
emellanåt	once in a while	0	0	1	0
emellanåt	occasionally	0	0	1	1
fontsizes	fontsizes	0	0	1	0
förbjöd	forbade	0	0	1	0
förbjöd	forbid	0	0	1	0
kapitalistiska	capitalistic	0	0	1	0
kapitalistiska	capitalist	0	0	1	0
sundsvall	sundsvall	0	0	1	0
kanadas	canada's	0	0	1	0
publicera	publish	0	0	1	1
abstrakta	abstract	0	0	1	0
talets	the speechs	0	0	1	0
talets	adding an s to the year.	0	0	1	0
talets	it means "decade" but would translate as "1950s"	0	0	1	0
talets	century	0	0	1	0
klitoris	clitoris	0	0	1	1
konstitutionen	constitution	0	0	1	0
förändrade	changed	0	0	1	0
förändrade	altered	0	0	1	0
tusen	thousands	0	0	1	0
tidskrifter	periodicals	0	0	1	0
tidskrifter	magazines	0	0	1	0
risk	risk	0	0	1	1
hörn	corner	0	0	1	1
ipredlagen	ipred act	0	0	1	0
satt	saat	0	0	1	0
satt	sat	0	0	1	0
nobelstiftelsen	nobel foundation	0	0	1	0
bonaparte	bonaparte	0	0	1	0
vintrar	winters	0	0	1	0
höra	hear	0	0	1	1
höra	know	0	0	1	0
höra	whore	0	0	1	0
begrepp	term	0	0	1	0
begrepp	concept	0	0	1	1
stöder	supporting	0	0	1	0
stöder	supports	0	0	1	0
armé	poor	0	0	1	0
armé	army	0	0	1	0
polis	police	0	0	1	1
autonoma	autonomous	0	0	1	0
autonoma	autonomic	0	0	1	0
sträng	string	0	0	1	1
sträng	strang	0	0	1	0
stilla	still	0	0	1	1
stilla	stationary	0	0	1	0
tycktes	tycktes	0	0	1	0
tycktes	seemed	0	0	1	0
hörs	heard	0	0	1	0
dödades	killed	0	0	1	0
dödades	were killed	0	0	1	0
värme	heat	0	0	1	1
värme	thermal	0	0	1	0
orsakar	causes	0	0	1	0
orsakas	caused	0	0	1	0
orsakas	causes	0	0	1	0
orsakas	caused by	0	0	1	0
orsakat	caused	0	0	1	0
utomeuropeiska	overseas	0	0	1	0
utomeuropeiska	non-european	0	0	1	0
startade	started	0	0	1	0
klarar	do	0	0	1	0
klarar	handle	0	0	1	0
president	president	0	0	1	1
orsakad	caused	0	0	1	0
orsakad	induced	0	0	1	0
indelat	divided	0	0	1	0
indelat	split	0	0	1	0
pågår	pagar	0	0	1	0
pågår	(in) progress	0	0	1	0
pågår	underway	0	0	1	0
indelas	divided	0	0	1	0
indelas	categorized	0	0	1	0
försök	experiments	0	0	1	0
försök	attempt	0	0	1	1
försök	expirements	0	0	1	0
höglandet	highlands	0	0	1	0
höglandet	the highland	0	0	1	0
bosättare	settlers	0	0	1	0
längsta	maximum	0	0	1	0
längsta	longest	0	0	1	0
indisk	indian	0	0	1	1
kvicksilver	mercury	0	0	1	1
kvicksilver	quicksilver	0	0	1	1
kvicksilver	witty zeal	0	0	1	0
fifa	fifa	0	0	1	0
panthera	panthera	0	0	1	0
belgien	belgium	0	0	1	1
munnen	the mouth	0	0	1	0
munnen	mouth	0	0	1	0
murray	murray	0	0	1	0
helena	helena	0	0	1	0
buddhister	budhists	0	0	1	0
buddhister	buddhists	0	0	1	0
arbetsgivaren	employer	0	0	1	0
besök	visit	0	0	1	1
nationell	national	0	0	1	1
personal	personal	0	0	1	0
personal	employed	0	0	1	0
personal	staff	0	0	1	1
rekord	record	0	0	1	1
amerikanen	american	0	0	1	0
amerikanen	the american	0	0	1	0
amerikaner	american	0	0	1	0
amerikaner	americans	0	0	1	0
irans	iran's	0	0	1	0
federationen	federation	0	0	1	0
federationen	the federation	0	0	1	0
gått	gone	0	0	1	0
gått	passed	0	0	1	0
friska	healthy	0	0	1	0
friska	fresh	0	0	1	0
friska	healty	0	0	1	0
aborter	abortions	0	0	1	0
infektioner	infections	0	0	1	0
infektioner	infection	0	0	1	0
aston	undra	0	0	1	0
aston	aston	0	0	1	0
aston	överraska	0	0	1	0
startat	started	0	0	1	0
medlemmar	members	0	0	1	0
förstörelse	destruction	0	0	1	1
downs	down	0	0	1	0
stimulerar	stimulates	0	0	1	0
stimulerar	stimulating	0	0	1	0
könsorgan	was organ	0	0	1	0
könsorgan	sex organ	0	0	1	0
könsorgan	genitals	0	0	1	1
miljon	one million	0	0	1	0
miljon	million	0	0	1	1
flamländska	flemish	0	0	1	0
myntades	coined	0	0	1	0
myntades	was coined	0	0	1	0
spåret	spparet	0	0	1	0
spåret	groove	0	0	1	0
spåret	track is	0	0	1	0
exakta	exact	0	0	1	0
huvudrollen	the main role	0	0	1	0
huvudrollen	leading part	0	0	1	0
listor	lists	0	0	1	0
luxemburg	luxemburg	0	0	1	0
luxemburg	luxembourg	0	0	1	1
tillvaron	existence	0	0	1	0
tillvaron	life	0	0	1	0
tillvaron	the subsistence	0	0	1	0
sida	website	0	0	1	0
sida	page	0	0	1	1
sida	side	0	0	1	1
side	side	0	0	1	0
kammaren	chamber	0	0	1	0
kammaren	the chamber	0	0	1	0
spåren	the tracks	0	0	1	0
spåren	tracks	0	0	1	0
spåren	wake	0	0	1	0
lägret	the camp	0	0	1	0
lägret	camp	0	0	1	0
tillät	distillate	0	0	1	0
tillät	allowed	0	0	1	0
röka	smoking	0	0	1	0
röka	roka	0	0	1	0
röka	smoke	0	0	1	1
liga	compatible	0	0	1	0
liga	league	0	0	1	1
mediet	medium	0	0	1	0
mediet	the medium	0	0	1	0
medier	media	0	0	1	0
medier	medias	0	0	1	0
väpnade	armed	0	0	1	0
milan	milan	0	0	1	0
anhängare	followers	0	0	1	0
anhängare	supporters	0	0	1	0
aids	aids	0	0	1	1
fängslades	imprisoned; jailed	0	0	1	0
fängslades	jailed	0	0	1	0
fängslades	gaoled; incarcerated	0	0	1	0
kiev	kiev	0	0	1	0
uppsala	uppsala	0	0	1	0
talet	rate	0	0	1	0
talet	century	0	0	1	0
tjänstemän	officals	0	0	1	0
tjänstemän	officers of	0	0	1	0
tjänstemän	officials	0	0	1	0
linköpings	linkopingas	0	0	1	0
linköpings	linköpings	0	0	1	0
linköpings	linköping's	0	0	1	0
ihop	up	0	0	1	0
ihop	together	0	0	1	1
talen	rate	0	0	1	0
talen	years	0	0	1	0
sluta	stop	0	0	1	1
sluta	end	0	0	1	1
ordförande	chairman	0	0	1	1
lämnade	did	0	0	1	0
lämnade	left	0	0	1	0
bestod	was	0	0	1	0
foto	photo	0	0	1	1
neutroner	neutrons	0	0	1	0
neutroner	neutron	0	0	1	0
larssons	larsson's	0	0	1	0
normer	norms	0	0	1	0
normer	standards	0	0	1	0
nietzsche	nietzsche	0	0	1	0
nomineringar	nominations	0	0	1	0
övergång	transition	0	0	1	1
folkvalda	elected	0	0	1	0
folkvalda	popularly elected	0	0	1	0
faktum	fact	0	0	1	1
iso	iso	0	0	1	0
reinfeldt	reinfeld	0	0	1	0
reinfeldt	reinfeldt	0	0	1	0
representant	representative	0	0	1	1
avslöjar	reveals	0	0	1	0
avslöjar	avslojar	0	0	1	0
starta	start	0	0	1	1
starta	startup	0	0	1	0
starta	launch	0	0	1	1
stewart	stewart	0	0	1	0
revolutionära	revolutionary	0	0	1	0
tävling	competition	0	0	1	1
tävling	contest	0	0	1	1
jordanien	jordan	0	0	1	1
engelskspråkiga	english-speaking	0	0	1	0
engelskspråkiga	the english language	0	0	1	0
arrangeras	(is) arranged	0	0	1	0
arrangeras	arranged	0	0	1	0
arrangeras	arrange	0	0	1	0
skalvet	quake	0	0	1	0
leddes	passed	0	0	1	0
leddes	was led	0	0	1	0
massiv	massive	0	0	1	1
månen	the moon	0	0	1	0
månen	man	0	0	1	0
objektet	the object	0	0	1	0
objektet	object	0	0	1	0
girls	girls	0	0	1	0
vikingatiden	the viking age	0	0	1	0
vikingatiden	vikings	0	0	1	0
omgående	immediately	0	0	1	1
omgående	immediate	0	0	1	1
objekten	items	0	0	1	0
objekten	objects	0	0	1	0
objekten	the objects	0	0	1	0
hollywood	hollywood	0	0	1	0
markerar	selects	0	0	1	0
markerar	marks	0	0	1	0
göras	made	0	0	1	0
göras	be made	0	0	1	0
göras	be made through	0	0	1	0
medeltiden	middle ages	0	0	1	0
besegrades	defeated	0	0	1	0
skaffade	acquired	0	0	1	0
skaffade	aquired	0	0	1	0
skaffade	took	0	0	1	0
sabbath	sabbath	0	0	1	0
göran	göran	0	0	1	0
göran	request	0	0	1	0
symptom	symptoms	0	0	1	0
symptom	symptom	0	0	1	1
hundar	dogs	0	0	1	0
götaland	götaland	0	0	1	0
götaland	gotaland	0	0	1	0
formell	formal	0	0	1	1
kontrast	contrast	0	0	1	1
möjliggjorde	made possible	0	0	1	0
möjliggjorde	enabled	0	0	1	0
möjliggjorde	allowed	0	0	1	0
troligtvis	probably	0	0	1	1
rådgivare	counsellor	0	0	1	1
rådgivare	advisor	0	0	1	1
östasien	east asia	0	0	1	0
bobo	bobo	0	0	1	0
palace	palace	0	0	1	0
stadsdelen	the district	0	0	1	0
stadsdelen	district	0	0	1	0
mina	my	0	0	1	0
mina	mine	0	0	1	1
modern	modern	0	0	1	1
mind	mind	0	0	1	0
triangel	triangle	0	0	1	1
drömmar	dreams	0	0	1	0
kolväten	hydrocarbons	0	0	1	0
kolväten	the hydrocarbon	0	0	1	0
skildringar	scenes	0	0	1	0
skildringar	description	0	0	1	0
skildringar	descriptions	0	0	1	0
tidiga	early	0	0	1	0
blåvitt	bluewhite	0	0	1	0
blåvitt	blåvitt	0	0	1	0
blåvitt	blue and white	0	0	1	0
europarådet	council of europe	0	0	1	0
europarådet	european council	0	0	1	0
muskler	muscles	0	0	1	0
bakgrunden	background	0	0	1	0
ulrich	ulrich	0	0	1	0
ep	ep	0	0	1	0
blue	blue	0	0	1	0
dessa	this	0	0	1	0
dessa	these	0	0	1	1
bildar	serves as	0	0	1	0
bildar	form	0	0	1	0
bildas	formed; made up (of)	0	0	1	0
bildas	formed	0	0	1	0
norra	north	0	0	1	1
norra	northern	0	0	1	1
inbördeskriget	civil war; civil war	0	0	1	0
inbördeskriget	civil war	0	0	1	0
godkänt	approved	0	0	1	0
godkänt	pass	0	0	1	0
påsken	easter	0	0	1	0
mario	mario	0	0	1	0
efterträdare	successor	0	0	1	1
luthers	luthers	0	0	1	0
luthers	luther's	0	0	1	0
luthers	luther	0	0	1	0
marie	marie	0	0	1	0
typ	kind of	0	0	1	0
typ	type	0	0	1	1
diskuterats	been discussed	0	0	1	0
diskuterats	discussed	0	0	1	0
maria	maria	0	0	1	0
don	don	0	0	1	1
dom	judgement	0	0	1	1
dom	conviction	0	0	1	0
materiella	material	0	0	1	0
talanger	talents	0	0	1	0
dog	died	0	0	1	0
slipknot	slipknot	0	0	1	0
stjärnan	star	0	0	1	0
stjärnan	the star	0	0	1	0
points	point	0	0	1	0
dos	dosage	0	0	1	1
dop	baptismal	0	0	1	0
dop	baptism	0	0	1	1
uttalande	statement	0	0	1	0
kristen	christian	0	0	1	1
feminister	feminists	0	0	1	0
koppla	coupling	0	0	1	0
koppla	connect	0	0	1	1
utom	except	0	0	1	1
utom	out	0	0	1	0
sjöfarten	maritime transport	0	0	1	0
sjöfarten	shipping	0	0	1	0
kronprins	crown prince	0	0	1	1
liza	liza	0	0	1	0
droger	drugs	0	0	1	0
skyldig	responsible	0	0	1	0
skyldig	guilty	0	0	1	1
slår	states	0	0	1	0
slår	switch	0	0	1	0
slår	beats	0	0	1	0
slås	beat	0	0	1	0
slås	is hit	0	0	1	0
slås	slas	0	0	1	0
bidrag	contribution	0	0	1	1
bidrag	contributions	0	0	1	0
odling	cultivation	0	0	1	1
utmärks	are characterized	0	0	1	0
utmärks	characterized	0	0	1	0
utmärkt	excellently	0	0	1	0
utmärkt	excellent; superb; marked by; characterized by	0	0	1	0
utmärkt	excellent	0	0	1	0
folke	folke	0	0	1	0
helhet	entirety	0	0	1	1
helhet	whole	0	0	1	1
vätet	hydrogen	0	0	1	0
vätet	the hydrogen	0	0	1	0
monica	monica	0	0	1	0
stycke	piece	0	0	1	1
stycke	piece; part; section	0	0	1	0
födelsetal	birthrate	0	0	1	1
födelsetal	birth rate	0	0	1	0
gällde	applied	0	0	1	0
gällde	was	0	0	1	0
gällde	applied to	0	0	1	0
ända	as far as	0	0	1	0
ända	up	0	0	1	0
meningar	sentences	0	0	1	0
dramaten	dramaten	0	0	1	0
stop	stop	0	0	1	0
vädret	weather	0	0	1	0
vädret	the weather	0	0	1	0
stor	big; great	0	0	1	0
stor	large	0	0	1	1
stor	great	0	0	1	1
stol	chair	0	0	1	1
stol	seat	0	0	1	1
strategiska	strategical	0	0	1	0
strategiska	strategic	0	0	1	0
christopher	christopher	0	0	1	0
stod	stood	0	0	1	0
earl	earl	0	0	1	0
bar	bar	0	0	1	1
bas	base	0	0	1	1
existerar	exists	0	0	1	0
skrivas	written	0	0	1	0
skrivas	printed	0	0	1	0
inlett	started	0	0	1	0
inlett	ushered in	0	0	1	0
inlett	initiated	0	0	1	0
existerat	existed	0	0	1	0
anlades	founded	0	0	1	0
anlades	were built	0	0	1	0
anlades	was built	0	0	1	0
bad	bath	0	0	1	1
fokus	focus	0	0	1	1
liggande	placed	0	0	1	0
liggande	overhead	0	0	1	0
liggande	lie	0	0	1	0
anknytning	tie	0	0	1	0
anknytning	link	0	0	1	0
anknytning	related	0	0	1	0
sänka	lower	0	0	1	1
sänka	marshy	0	0	1	0
förlag	publishers	0	0	1	0
förlag	magazine	0	0	1	0
förlag	forlag	0	0	1	0
avvikande	different	0	0	1	0
avvikande	deviant; divergent; different	0	0	1	0
zonen	the zone	0	0	1	0
zonen	zone	0	0	1	0
zoner	zones	0	0	1	0
gunnar	gunnar	0	0	1	0
dittills	thus far	0	0	1	0
dittills	so far	0	0	1	0
växer	growing	0	0	1	0
växer	grows	0	0	1	0
inledningsvis	initially	0	0	1	0
inledningsvis	in the beginning	0	0	1	0
inledningsvis	by way of introduction	0	0	1	1
avgörs	determined	0	0	1	0
avgörs	is determined	0	0	1	0
avgörs	decided	0	0	1	0
skrevs	written	0	0	1	0
skrevs	was	0	0	1	0
hergé	herge	0	0	1	0
hergé	hergé	0	0	1	0
naturligtvis	course	0	0	1	0
naturligtvis	off course	0	0	1	0
naturligtvis	naturally	0	0	1	1
skrift	no.	0	0	1	0
skrift	book	0	0	1	0
skrift	writing	0	0	1	1
oförmåga	inability	0	0	1	1
oförmåga	failure	0	0	1	0
oförmåga	incapacity	0	0	1	1
sorts	variety	0	0	1	0
omkringliggande	surrounding	0	0	1	0
omkringliggande	neighbouring	0	0	1	0
avgöra	decide	0	0	1	1
avgöra	determine	0	0	1	1
smguld	swedish championship gold	0	0	1	0
smguld	gold medal in the swedish championships	0	0	1	0
smguld	sm gold	0	0	1	0
artikel	article	0	0	1	1
örebro	Örebro	0	0	1	0
jämförelsevis	comparative	0	0	1	0
jämförelsevis	in comparison	0	0	1	0
jämförelsevis	comparatively	0	0	1	1
armeniska	armenian	0	0	1	0
nationalister	nationalists	0	0	1	0
innehåll	content	0	0	1	1
innehåll	contents	0	0	1	1
motto	motto	0	0	1	1
behöver	need	0	0	1	0
förhöjd	elevated	0	0	1	0
förhöjd	enhanced	0	0	1	0
regelbundet	regularly	0	0	1	1
regelbundet	regularily	0	0	1	0
isotoper	isotopes	0	0	1	0
fns	un's	0	0	1	0
fns	tris	0	0	1	0
regering	the government	0	0	1	0
regering	government	0	0	1	1
und	und	0	0	1	0
ung	young	0	0	1	1
ernst	ernst	0	0	1	0
regelbunden	regular	0	0	1	1
obamas	obama's	0	0	1	0
obamas	obamas	0	0	1	0
obamas	obama	0	0	1	0
uno	uno	0	0	1	0
mellanrum	gap	0	0	1	1
mellanrum	space	0	0	1	1
hjärna	brain	0	0	1	1
föregångare	predecessor	0	0	1	0
föregångare	precursor	0	0	1	1
sägas	is said	0	0	1	0
sägas	is said (to be)	0	0	1	0
sägas	said	0	0	1	0
flickvän	girlfriend	0	0	1	1
avsikt	intention	0	0	1	1
avsikt	intends	0	0	1	0
sommartid	summer-time	0	0	1	0
sommartid	summer	0	0	1	0
sommartid	during summer	0	0	1	0
mördades	murdered	0	0	1	0
mördades	was murdered	0	0	1	0
mördades	murder was	0	0	1	0
studerar	study	0	0	1	0
studerar	studies	0	0	1	0
omstritt	controversial	0	0	1	0
varmt	hot	0	0	1	0
varmt	warm	0	0	1	0
basis	basis	0	0	1	1
studerat	studied	0	0	1	0
blodkroppar	blood cells	0	0	1	0
blodkroppar	corpuscle	0	0	1	0
cyrus	cyrus	0	0	1	0
ting	things	0	0	1	0
ting	matters	0	0	1	0
ting	thing	0	0	1	1
frisk	healthy	0	0	1	1
frisk	fresh	0	0	1	1
åtal	prosecution	0	0	1	1
idol	idol	0	0	1	1
minoriteten	minority	0	0	1	0
betydelsefull	meningful	0	0	1	0
betydelsefull	significant	0	0	1	1
förhållandet	the ratio	0	0	1	0
förhållandet	the relation	0	0	1	0
förhållandet	relationship	0	0	1	0
provinsen	province	0	0	1	0
provinsen	rovisen	0	0	1	0
provinsen	the province	0	0	1	0
utseende	appearance	0	0	1	1
förhållanden	relationships	0	0	1	0
förhållanden	conditions	0	0	1	0
förhållanden	n/a	0	0	1	0
mindre	smaller	0	0	1	1
mindre	less	0	0	1	1
hårt	hard	0	0	1	1
hårt	resin	0	0	1	0
hårt	difficult	0	0	1	0
etniskt	ethnical	0	0	1	0
etniskt	ethnic	0	0	1	0
azerbajdzjan	azerbaijan	0	0	1	0
azerbajdzjan	azerbaijani	0	0	1	0
say	say	0	0	1	0
angående	concerning	0	0	1	1
angående	reference	0	0	1	0
etniska	ethnic	0	0	1	0
tillhörighet	affiliation	0	0	1	0
tillhörighet	belonging	0	0	1	1
tillhörighet	belonging; affiliation	0	0	1	0
ära	oar	0	0	1	0
ära	glory	0	0	1	1
ära	honor	0	0	1	1
pornografi	pornography	0	0	1	1
paradiset	the paradise	0	0	1	0
paradiset	paradise	0	0	1	0
ix	4	0	0	1	0
ix	the ninth	0	0	1	0
albaner	albanians	0	0	1	0
mexico	mexico	0	0	1	1
kvinnor	female	0	0	1	0
kvinnor	women	0	0	1	1
ip	ip	0	0	1	0
sushi	sushi	0	0	1	0
iu	iu	0	0	1	0
it	it	0	0	1	0
benämningar	terms	0	0	1	0
benämningar	names	0	0	1	0
ii	(ii)	0	0	1	0
cant	cant	0	0	1	0
dokument	files	0	0	1	0
dokument	document	0	0	1	1
dokument	documents	0	0	1	0
im	im	0	0	1	0
il	il	0	0	1	0
jesu	jesus	0	0	1	0
jesu	jesu	0	0	1	0
colosseum	colosseum	0	0	1	0
strömmen	current	0	0	1	0
strömmen	the stream	0	0	1	0
stoppa	stop	0	0	1	1
konkurrensen	the competition	0	0	1	0
konkurrensen	competitive	0	0	1	0
make	make	0	0	1	0
make	husband	0	0	1	1
redaktör	editor	0	0	1	1
bella	bella	0	0	1	0
kommunistpartiets	communist party	0	0	1	0
kommunistpartiets	the communist partys	0	0	1	0
kommunistpartiets	the communist party	0	0	1	0
roland	roland	0	0	1	0
industriell	industrial	0	0	1	1
makt	power	0	0	1	1
anglosaxiska	anglo-saxon	0	0	1	0
högtryck	anticyclone	1	1	0	0
högtryck	flat out	1	0	1	0
högtryck	the heat is on	1	0	1	0
högtryck	hotryck	1	0	1	0
högtryck	high pressure	1	0	1	1
högtryck	pressure	1	0	1	0
högtryck	high presssure	1	0	1	0
högtryck	he	1	0	1	0
dillinger	dillinger	0	0	1	0
explosionen	the explosion	0	0	1	0
kim	kim	0	0	1	0
nicklas	niclas	0	0	1	0
nicklas	nicklas	0	0	1	0
folkrikaste	populous	0	0	1	0
folkrikaste	people rich	0	0	1	0
folkrikaste	most populus	0	0	1	0
akademiska	academical	0	0	1	0
akademiska	academic	0	0	1	0
protesterna	protests	0	0	1	0
protesterna	the protests	0	0	1	0
roms	rome's	0	0	1	0
roms	roms	0	0	1	0
roms	romes	0	0	1	0
vetenskaplig	learn scientific	0	0	1	0
vetenskaplig	scientific	0	0	1	1
sydamerika	south america	0	0	1	1
städer	urban	0	0	1	0
städer	cities	0	0	1	0
roma	roma	0	0	1	0
slå	beat	0	0	1	1
slå	hit	0	0	1	1
slå	sla	0	0	1	0
viktiga	important	0	0	1	0
facto	facto	0	0	1	0
just	right	0	0	1	1
just	currently	0	0	1	0
just	just	0	0	1	1
diameter	diameter	0	0	1	1
sporting	sporting	0	0	1	0
universitet	university	0	0	1	1
psykos	phychosis	0	0	1	0
psykos	psychosis	0	0	1	1
bollen	the ball	0	0	1	0
bollen	ball	0	0	1	0
styrelsen	the board	0	0	1	0
styrelsen	board	0	0	1	0
human	human	0	0	1	0
anders	anders	0	0	1	0
beskriver	describes	0	0	1	0
fysiker	physicist	0	0	1	1
fysiker	physicists	0	0	1	0
skulptur	sculpture	0	0	1	1
troligt	likely	0	0	1	1
royal	royal	0	0	1	0
julen	julien	0	0	1	0
julen	christmas	0	0	1	0
memoarer	memoirs	0	0	1	1
jules	jules	0	0	1	0
friedrich	friedrich	0	0	1	0
ökat	increased	0	0	1	0
amerikas	america	0	0	1	0
amerikas	america's	0	0	1	0
harald	harald	0	0	1	0
borgen	castle	0	0	1	0
borgen	bail	0	0	1	1
borgen	the castle	0	0	1	0
komintern	comintern	0	0	1	0
komintern	komintern	0	0	1	0
arkitekturen	the architecture	0	0	1	0
arkitekturen	architecture	0	0	1	0
gustav	gustav	0	0	1	0
typiskt	typically	0	0	1	1
typiskt	typical	0	0	1	0
utrikesminister	minister of foreign affairs	0	0	1	0
utrikesminister	foreign minister	0	0	1	0
tittar	looking; viewing; viewer	0	0	1	0
tittar	viewing	0	0	1	0
lösning	solution	0	0	1	1
lösning	solution; resolution	0	0	1	0
gustaf	gustaf	0	0	1	0
trafikeras	served	0	0	1	0
trafikeras	trafficked	0	0	1	0
trafikerar	traffic	0	0	1	0
trafikerar	frequent	0	0	1	0
västerbottens	västerbottens	0	0	1	0
västerbottens	west bothnia	0	0	1	0
västerbottens	västerbotten's	0	0	1	0
medborgarskap	citizenship	0	0	1	1
kommunerna	kommunera	0	0	1	0
kommunerna	municipalities	0	0	1	0
kommunerna	the municipalities	0	0	1	0
intensiv	intensity	0	0	1	0
intensiv	intense	0	0	1	1
litauen	lithuania	0	0	1	1
syrien	syria	0	0	1	1
kemiska	chemical	0	0	1	0
vattnet	water	0	0	1	0
vattnet	the water	0	0	1	0
kontinent	continent	0	0	1	1
kunna	to	0	0	1	0
kunna	be able	0	0	1	0
eker	spoke	1	1	0	1
dead	dead	0	0	1	0
pär	pär	0	0	1	0
befolkningen	the population	0	0	1	0
befolkningen	population	0	0	1	0
förklaringar	explanations	0	0	1	0
jupiter	jupiter	0	0	1	1
befann	found	0	0	1	0
befann	located	0	0	1	0
kemiskt	chemically	0	0	1	0
dominerade	dominated	0	0	1	0
tappar	drop	0	0	1	0
tappar	lose	0	0	1	0
statistik	statistics	0	0	1	1
oralsex	oral sex	0	0	1	0
teoretiska	theoretical	0	0	1	0
nervosa	nervosa	0	0	1	0
shakespeare	shakespeare	0	0	1	0
gåva	gift	0	0	1	1
filmatiserats	cinematized	0	0	1	0
filmatiserats	been filmed	0	0	1	0
filmatiserats	screened	0	0	1	0
dödshjälp	euthanasy	0	0	1	0
dödshjälp	euthanasia	0	0	1	1
knep	tricks	0	0	1	0
knep	sleight of hand	0	0	1	0
angrepp	attack	0	0	1	1
grannländerna	neighbors	0	0	1	0
grannländerna	neighbouring countries	0	0	1	0
burj	burj	0	0	1	0
versioner	versions	0	0	1	0
bolt	bolt	0	0	1	0
burr	burr	0	0	1	0
stjärna	star	0	0	1	1
super	super	0	0	1	0
naturtillgångar	natural resources	0	0	1	0
flyttat	moved	0	0	1	0
maskiner	equipment	0	0	1	0
maskiner	machines	0	0	1	0
teoretiskt	theoretic	0	0	1	0
teoretiskt	theoretical	0	0	1	0
mycket	very	0	0	1	1
mycket	much	0	0	1	1
tillverkar	makes	0	0	1	0
tillverkar	producing	0	0	1	0
tillverkar	manufactures	0	0	1	0
tillverkas	is made	0	0	1	0
tillverkas	manufacture	0	0	1	0
tillverkas	manufactured	0	0	1	0
magazine	magazine	0	0	1	0
ishockey	ice hockey	0	0	1	1
ishockey	hockey	0	0	1	0
grenen	the branch	0	0	1	0
grenen	branch	0	0	1	0
psykisk	psychic	0	0	1	1
psykisk	mental	0	0	1	0
romantiska	romantic	0	0	1	0
verkställande	executive	0	0	1	1
jens	jens	0	0	1	0
poäng	score	0	0	1	0
poäng	point	0	0	1	1
romulus	romulus	0	0	1	0
orsak	reason	0	0	1	1
orsak	cause	0	0	1	1
orsak	factor	0	0	1	0
down	down	0	0	1	0
utbildning	education	0	0	1	1
utbildning	eduction	0	0	1	0
utbildning	education and training	0	0	1	0
amsterdam	amsterdam	0	0	1	0
svartån	svartån	0	0	1	0
svartån	svartån (black stream)	0	0	1	0
fastlandet	mainland	0	0	1	0
platån	sycamore	0	0	1	0
platån	the plateau	0	0	1	0
platån	plateau	0	0	1	0
estniska	estonian	0	0	1	1
tennis	tennis	0	0	1	1
rådets	council	0	0	1	0
närheten	near	0	0	1	0
närheten	the vicinity	0	0	1	0
bolivia	bolivia	0	0	1	1
över	of	0	0	1	1
över	over	0	0	1	1
påföljande	following	0	0	1	1
påföljande	subsequent	0	0	1	1
hyllade	celebrated	0	0	1	0
hyllade	acclaimed	0	0	1	0
form	form	0	0	1	1
präglad	characterize	0	0	1	0
präglad	characterized	0	0	1	0
präglad	marked	0	0	1	0
norrlands	northern sweden's	0	0	1	0
norrlands	lapland's	0	0	1	0
norrlands	norrland	0	0	1	0
batman	batman	0	0	1	0
ford	ford	0	0	1	0
präglas	characterised	0	0	1	0
präglas	characterized	0	0	1	0
återstår	remains	0	0	1	0
återstår	remain	0	0	1	0
berätta	tell	0	0	1	1
bero	depend	0	0	1	1
bero	due	0	0	1	0
byggde	was	0	0	1	0
byggde	founded (on)	0	0	1	0
byggde	built	0	0	1	0
definierade	defined	0	0	1	0
tempel	temple	0	0	1	1
spelade	played	0	0	1	0
långvarig	of long duration	0	0	1	0
långvarig	prolonged; lengthy; long	0	0	1	0
långvarig	long	0	0	1	1
hjälper	helps	0	0	1	0
hjälper	shows	0	0	1	0
positiv	positive	0	0	1	1
slaviska	slav	0	0	1	0
slaviska	slavic	0	0	1	1
slaviska	slavonic	0	0	1	1
bränsle	fuel	0	0	1	1
flygande	flying	0	0	1	1
skelett	skeleton	0	0	1	1
beteckningen	the label	0	0	1	0
beteckningen	designation.........	0	0	1	0
beteckningen	designation	0	0	1	0
avsnitt	section	0	0	1	1
avsnitt	part	0	0	1	1
avsnitt	episode	0	0	1	1
frihetliga	libertarian	0	0	1	0
förnuft	common sense	0	0	1	0
förnuft	reason	0	0	1	1
skåne	skåne	0	0	1	0
skåne	scania	0	0	1	1
välkända	known	0	0	1	0
välkända	well known	0	0	1	0
socialdemokrater	social democrats	0	0	1	0
uttryckligen	explicitly	0	0	1	0
uttryckligen	specifically	0	0	1	0
spänningen	exitement	0	0	1	0
spänningen	voltage	0	0	1	0
handelspartner	trading partner	0	0	1	0
tosh	tosh	0	0	1	0
kanske	may	0	0	1	0
världskrigets	the world war's	0	0	1	0
världskrigets	world war	0	0	1	0
månaderna	months	0	0	1	0
månaderna	are compelled	0	0	1	0
många	many	0	0	1	1
långsammare	more slowly	0	0	1	0
långsammare	slower	0	0	1	0
primtal	prime number	0	0	1	0
byggnaden	building	0	0	1	0
byggnaden	the building	0	0	1	0
vista	vista	0	0	1	0
handen	the hand	0	0	1	0
handen	hand	0	0	1	0
handel	commercial	0	0	1	0
handel	trade	0	0	1	1
kunnat	could	0	0	1	0
kunnat	could have been	0	0	1	0
kunnat	been	0	0	1	0
betala	pay	0	0	1	1
följaktligen	consequently	0	0	1	1
digital	digital	0	0	1	1
betalt	charge	0	0	1	0
marxism	marxism	0	0	1	0
kungamakten	monarchy	0	0	1	0
kungamakten	the monarchy	0	0	1	0
lågt	low	0	0	1	1
löpande	running	0	0	1	0
löpande	assembly	0	0	1	0
löpande	conveyor (belt)	0	0	1	0
stöter	thrust	0	0	1	0
stöter	run	0	0	1	0
frodo	frodo	0	0	1	0
exporten	exports	0	0	1	0
exporten	the export	0	0	1	0
jones	jones	0	0	1	0
drivs	driven	0	0	1	0
drivs	run	0	0	1	0
drivs	powered	0	0	1	0
accepterade	accepted	0	0	1	0
salt	salt	0	0	1	1
riktad	directed	0	0	1	0
frigörelse	liberation	0	0	1	1
fss	fss	0	0	1	0
expandera	expand	0	0	1	1
undervisade	taught	0	0	1	0
riktat	riktag	0	0	1	0
riktat	directed	0	0	1	0
riktat	pointed	0	0	1	0
riktas	directed (at)	0	0	1	0
riktas	direct	0	0	1	0
riktas	target	0	0	1	0
riktar	targets	0	0	1	0
riktar	target	0	0	1	0
milt	mild	0	0	1	0
armar	arms	0	0	1	0
bomben	bomb	0	0	1	0
bomben	the bomb	0	0	1	0
telefon	telephone	0	0	1	1
sanna	true	0	0	1	0
mild	mild	0	0	1	1
mild	soft	0	0	1	1
bomber	bombs	0	0	1	0
blåser	blows	0	0	1	0
blåser	blowing	0	0	1	0
vikingarna	the vikings	0	0	1	0
stulna	stolen	0	0	1	0
människan	the human	0	0	1	0
människan	people	0	0	1	0
människan	man	0	0	1	0
imperiet	the empire	0	0	1	0
imperiet	empire	0	0	1	0
beträffande	on	0	0	1	0
avbrott	break	0	0	1	1
avbrott	breaks	0	0	1	0
uppdelning	division	0	0	1	1
uppdelning	partitioning	0	0	1	0
uppdelning	playback	0	0	1	0
reptiler	reptiles	0	0	1	0
människas	human's; man's	0	0	1	0
människas	human	0	0	1	0
byggnadsverk	building	0	0	1	0
byggnadsverk	construction	0	0	1	0
byggnadsverk	edifice	0	0	1	0
me	me	0	0	1	0
farlig	dangerous	0	0	1	1
farlig	hazardous	0	0	1	1
skapad	created	0	0	1	0
vetenskapsmän	scientist	0	0	1	0
vetenskapsmän	scientists	0	0	1	0
illa	bad	0	0	1	0
hösten	the autumn	0	0	1	0
hösten	the fall	0	0	1	0
hösten	fall	0	0	1	0
din	yours	0	0	1	1
din	your	0	0	1	1
apartheid	apartheid	0	0	1	1
dig	up	0	0	1	0
trenden	trend	0	0	1	0
trenden	the trend	0	0	1	0
kupol	regularly	1	0	1	0
kupol	cupola	1	1	0	1
kupol	dome	1	1	0	1
kupol	regular	1	0	1	0
kupol	combatant	1	0	1	0
kupol	cu	1	0	1	0
afrikansk	african	0	0	1	1
dit	there	0	0	1	1
dit	where	0	0	1	1
tillräcklig	sufficient	0	0	1	1
tillräcklig	enough	0	0	1	1
bulgarien	bulgaria	0	0	1	1
olympia	olympia	0	0	1	0
ville	wanted (to)	0	0	1	0
ville	did	0	0	1	0
ville	wanted	0	0	1	0
diskografi	discography	0	0	1	0
villa	house	0	0	1	0
villa	villa	0	0	1	1
slagit	held	0	0	1	0
slagit	beaten	0	0	1	0
reklamen	the commercial	0	0	1	0
reklamen	commercial; ad; advertisment	0	0	1	0
reklamen	advertising	0	0	1	0
invandringen	immigration	0	0	1	0
ökande	increasing	0	0	1	1
ökande	rising	0	0	1	0
rymden	space	0	0	1	0
uppväxt	growing up	0	0	1	0
fäste	bracket	0	0	1	0
fäste	attachment	0	0	1	1
bakom	behind	0	0	1	1
högra	right	0	0	1	0
kännedom	known	0	0	1	0
kännedom	knowledge	0	0	1	1
högre	higher	0	0	1	1
vanligen	usually	0	0	1	1
vanligen	typically	0	0	1	0
afghanistan	afghanisthan	0	0	1	0
afghanistan	afghanistan	0	0	1	1
varpå	thereafter	0	0	1	0
varpå	whereupon	0	0	1	1
varpå	after which	0	0	1	0
viktig	major	0	0	1	0
viktig	important	0	0	1	1
kokain	cocaine	0	0	1	1
kokain	cocain	0	0	1	0
kompositörer	composers	0	0	1	0
kompositörer	compositors	0	0	1	0
bibliotek	library	0	0	1	1
lennon	lennon	0	0	1	0
bekämpa	prevent	0	0	1	0
bekämpa	combat; fight	0	0	1	0
bekämpa	fight	0	0	1	1
international	international	0	0	1	1
avsluta	finish	0	0	1	1
avsluta	exit	0	0	1	0
nationalismen	nationalism	0	0	1	0
tibet	tibet	0	0	1	0
mr	herr	0	0	1	0
mr	mr	0	0	1	0
utlänningar	foreigners	0	0	1	0
avsaknad	absence	0	0	1	0
specialiserade	specialized	0	0	1	0
specialiserade	special	0	0	1	0
kommun	local	0	0	1	0
kommun	municipality	0	0	1	1
beskrivits	described	0	0	1	0
boy	boy	0	0	1	0
diagnoser	diagnoses	0	0	1	0
canadian	canadian	0	0	1	0
institute	institute	0	0	1	0
bor	lives	0	0	1	0
gyllene	golden	0	0	1	1
gyllene	golden; gilded	0	0	1	0
folkmun	popular lore; popularly	0	0	1	0
folkmun	common speech	0	0	1	0
folkmun	colloquially	0	0	1	0
bok	book	0	0	1	1
bon	nests	0	0	1	0
bon	bon	0	0	1	0
extrem	extreme	0	0	1	1
bob	bob	0	0	1	0
nyfödda	newborn	0	0	1	0
bolivianska	bolivian	0	0	1	0
förbinder	connects	0	0	1	0
förbinder	undertake	0	0	1	0
departement	departement	0	0	1	0
departement	department	0	0	1	1
röstade	voted	0	0	1	0
ån	on	0	0	1	0
ån	from	0	0	1	0
ån	the river	0	0	1	0
dvärg	dwarf	0	0	1	1
sporter	sports	0	0	1	0
enorma	enormous	0	0	1	0
rösträtt	vote	0	0	1	0
rösträtt	right to vote	0	0	1	0
sporten	the sport	0	0	1	0
sporten	sport	0	0	1	0
sporten	port	0	0	1	0
religionsfrihet	freedom of religion	0	0	1	0
religionsfrihet	religious freedom	0	0	1	0
religionsfrihet	religion	0	0	1	0
åt	to	0	0	1	1
åt	for	0	0	1	1
ås	ridge	0	0	1	1
ås	site	0	0	1	0
år	the year	0	0	1	0
år	year	0	0	1	1
franco	franco	0	0	1	0
hemmaarena	home ground	0	0	1	0
hemmaarena	home field	0	0	1	0
tennisspelare	tennis player	0	0	1	0
socialister	socialists	0	0	1	0
semifinalen	the semi-final	0	0	1	0
semifinalen	semi finals	0	0	1	0
semifinalen	semifinal	0	0	1	0
särskilda	specific	0	0	1	0
särskilda	special	0	0	1	0
peru	peru	0	0	1	1
kristian	kristian	0	0	1	0
omöjligt	impossible	0	0	1	0
left|px	left px	0	0	1	0
ställdes	was positioned	0	0	1	0
ställdes	prepared	0	0	1	0
detaljer	details	0	0	1	0
avsattes	deposited	0	0	1	0
avsattes	dismissed	0	0	1	0
brukade	used to	0	0	1	0
brukade	used	0	0	1	0
kemisk	chemical	0	0	1	1
världsdel	continent	0	0	1	1
županija	country	0	0	1	0
snö	snow	0	0	1	1
fartyget	vessel	0	0	1	0
fartyget	ship; vessel	0	0	1	0
fartyget	boat	0	0	1	0
förknippad	associated	0	0	1	0
försäljning	sales	0	0	1	0
försäljning	sale	0	0	1	1
fly	escape	0	0	1	1
tokyo	tokyo	0	0	1	0
sångerna	song are	0	0	1	0
sångerna	the songs	0	0	1	0
soul	soul	0	0	1	0
kombination	combination	0	0	1	1
vittnen	witnesses	0	0	1	0
akademien	the academy	0	0	1	0
akademien	academy	0	0	1	0
akademien	riksdagens	0	0	1	0
anslutna	affiliated	0	0	1	0
anslutna	connected	0	0	1	0
bristande	lack of	0	0	1	0
bristande	lack	0	0	1	0
bristande	wanting	0	0	1	0
ulf	ulf	0	0	1	0
hiroshima	hiroshima	0	0	1	0
översättning	translation	0	0	1	1
översättning	translation thereof	0	0	1	0
kenneth	kenneth	0	0	1	0
uruguay	uruguay	0	0	1	0
erövringen	conquest	0	0	1	0
winston	winston	0	0	1	0
agent	agent	0	0	1	1
norrmän	norwegians	0	0	1	0
skadades	damaged	0	0	1	0
skadades	was wounded	0	0	1	0
council	council	0	0	1	0
asteroidbältet	asteroid belt	0	0	1	0
asteroidbältet	the asteroid belt	0	0	1	0
dennis	dennis	0	0	1	0
kunglig	royal	0	0	1	1
pink	pink	0	0	1	0
pink	piddle	0	0	1	1
erövring	conquest	0	0	1	1
diskuterades	discussed	0	0	1	0
oslo	oslo	0	0	1	1
varor	products	0	0	1	0
draperi	curtains	1	0	1	0
draperi	corresponding	1	0	1	0
draperi	acoording	1	0	1	0
draperi	drapery; curtain	1	0	1	0
draperi	daperi	1	1	0	0
draperi	curtian	1	1	0	0
draperi	curtain	1	1	0	1
draperi	drapery	1	1	0	1
ekonomiska	economic	0	0	1	0
ekonomiska	economical	0	0	1	0
till	to	0	0	1	1
årstiderna	seasons	0	0	1	0
årstiderna	the seasons	0	0	1	0
årstiderna	arstiderna	0	0	1	0
gitarrist	guitarist	0	0	1	1
nya	new	0	0	1	0
nya	severe	0	0	1	0
nye	new	0	0	1	0
mat	food	0	0	1	1
rökning	smoking	0	0	1	1
regeringstid	term of government	0	0	1	0
regeringstid	term of government; term of office	0	0	1	0
regeringstid	reign	0	0	1	0
may	may	0	0	1	0
thåström	thåström	0	0	1	0
thåström	thastrom	0	0	1	0
antogs	adoption	0	0	1	0
antogs	was assumed	0	0	1	0
centrum	center	0	0	1	1
maj	may	0	0	1	1
mao	mao	0	0	1	0
man	is	0	0	1	0
man	one	0	0	1	1
asien	asia	0	0	1	1
johnson	johnson	0	0	1	0
förekommit	occured	0	0	1	0
förekommit	occurred	0	0	1	0
q	q	0	0	1	0
tala	speaking	0	0	1	0
tala	speak	0	0	1	1
basket	basketball	0	0	1	0
romantiken	romance	0	0	1	0
romantiken	romanticism	0	0	1	0
undantag	exception	0	0	1	1
undantag	except	0	0	1	0
lsd	lsd	0	0	1	0
bussar	bus	0	0	1	0
bevisa	prove	0	0	1	1
alfabetet	alphabet	0	0	1	0
alfabetet	the alphabet	0	0	1	0
unionen	union	0	0	1	0
unionen	the union	0	0	1	0
unionen	european union	0	0	1	0
moralisk	moralic	0	0	1	0
moralisk	moral	0	0	1	1
huvudsak	in principal; chiefly	0	0	1	0
huvudsak	mainly	0	0	1	0
huvudsak	main thing	0	0	1	0
lyrik	poetry	0	0	1	0
group	group	0	0	1	0
landskap	province	0	0	1	1
landskap	landscapes	0	0	1	0
landskap	landscape	0	0	1	1
juryn	the selection panel	0	0	1	0
juryn	the jury	0	0	1	0
juryn	jury	0	0	1	0
dagbladet	daily paper	0	0	1	0
dagbladet	dagbladet	0	0	1	0
sekter	sects	0	0	1	0
inkomster	income	0	0	1	1
inkomster	revenue	0	0	1	0
rasen	breed	0	0	1	0
rasen	the race	0	0	1	0
policy	policy	0	0	1	0
main	main	0	0	1	0
texas	texas	0	0	1	0
steget	step	0	0	1	0
janeiro	janeiro	0	0	1	0
ibrahimović	ibrahimovic	0	0	1	0
förbättringar	improvements	0	0	1	0
förbättringar	improvement	0	0	1	0
stärkelse	starch	0	0	1	1
språkliga	linguistic	0	0	1	0
språkliga	language compatible	0	0	1	0
egenskaper	characteristics	0	0	1	0
egenskaper	charactiristics	0	0	1	0
egenskaper	qualities	0	0	1	0
sibirien	siberia	0	0	1	1
leds	led by	0	0	1	0
leds	passed	0	0	1	0
vindkraft	wind power	0	0	1	0
vindkraft	wind	0	0	1	0
uppskattning	appreciation	0	0	1	1
uppskattning	estimated	0	0	1	0
leda	lead	0	0	1	1
ledd	led	0	0	1	0
rock	rock	0	0	1	0
tysklands	germany's	0	0	1	0
tysklands	germanys	0	0	1	0
guevara	guevara	0	0	1	0
latin	latin	0	0	1	1
tacitus	tacitus	0	0	1	0
ännu	even	0	0	1	1
ännu	still	0	0	1	1
ännu	yet	0	0	1	1
sänts	sants	0	0	1	0
sänts	sent	0	0	1	0
hellre	rather	0	0	1	1
hellre	more preferably	0	0	1	0
ålder	age	0	0	1	1
ålder	alder	0	0	1	0
vattendrag	water	0	0	1	0
vattendrag	streams	0	0	1	0
vattendrag	watercourse	0	0	1	1
avkomma	progeny	0	0	1	1
avkomma	offspring	0	0	1	1
girl	girl	0	0	1	0
saudiarabien	saudi arabia	0	0	1	0
canada	canada	0	0	1	1
jackson	mrs. jackson	0	0	1	0
jackson	jackson	0	0	1	0
tillåtelse	allowed	0	0	1	0
tillåtelse	permission	0	0	1	1
pamela	pamela	0	0	1	0
hemmet	home	0	0	1	0
hemmet	the home	0	0	1	0
kattdjur	cat	0	0	1	1
kattdjur	felidae	0	0	1	0
kärnor	core	0	0	1	0
kärnor	cores	0	0	1	0
valdes	representatives'	0	0	1	0
valdes	selected	0	0	1	0
valdes	chosen; elected	0	0	1	0
rådande	current	0	0	1	1
rådande	prevalent	0	0	1	0
ansiktet	face	0	0	1	0
monster	monster	0	0	1	1
monster	monsters	0	0	1	0
ort	place	0	0	1	1
ort	neighborhood	0	0	1	0
ort	location	0	0	1	0
chiles	chiles	0	0	1	0
chiles	chile's	0	0	1	0
valrörelsen	election campaign	0	0	1	0
valrörelsen	the election campaign	0	0	1	0
oro	anxiety	0	0	1	1
oro	worry	0	0	1	1
oro	concern	0	0	1	1
ajax	ajax	0	0	1	0
california	california	0	0	1	0
brooke	brooke	0	0	1	0
kognitiva	cognitive	0	0	1	0
ord	word	0	0	1	1
ord	words	0	0	1	1
tunnelbanan	subway; tube; underground	0	0	1	0
tunnelbanan	the subway	0	0	1	0
tunnelbanan	metro	0	0	1	0
keith	keith	0	0	1	0
verkade	did	0	0	1	0
verkade	appeared to	0	0	1	0
verkade	worked	0	0	1	0
verkade	were active	0	0	1	0
verkade	was active	0	0	1	0
gott	good	0	0	1	1
gott	practically; good	0	0	1	0
anledning	reason	0	0	1	1
anledning	cause	0	0	1	1
preventivmedel	contraceptives	0	0	1	0
preventivmedel	preventivedel	0	0	1	0
östra	ostra	0	0	1	0
östra	eastern	0	0	1	1
våldet	the violence	0	0	1	0
våldet	violence	0	0	1	0
använts	was used	0	0	1	0
använts	used	0	0	1	0
uppvisar	shows	0	0	1	0
rankningar	ranking	0	0	1	0
rankningar	rankings	0	0	1	0
öde	fate	0	0	1	1
kraftig	strong	0	0	1	0
egentligen	actually	0	0	1	1
egentligen	actual	0	0	1	0
egentligen	really	0	0	1	1
first	first	0	0	1	0
centrala	central	0	0	1	0
grupperna	groups	0	0	1	0
intryck	impression	0	0	1	1
intryck	appearance	0	0	1	0
uttalanden	statements	0	0	1	0
rachel	rachel	0	0	1	0
folklig	popular	0	0	1	1
folklig	folk	0	0	1	0
biografen	the cinema	0	0	1	0
biografen	movie theater	0	0	1	0
biografen	cinema	0	0	1	0
centralt	central	0	0	1	0
centralt	centrally	0	0	1	0
skapandet	creation	0	0	1	0
skapandet	the making	0	0	1	0
kommunism	communism	0	0	1	1
mängden	amount	0	0	1	0
mängden	the amount	0	0	1	0
bronsåldern	bronze age	0	0	1	0
bronsåldern	the bronze age	0	0	1	0
grå	gray	0	0	1	1
grå	grey	0	0	1	1
alfred	alfred	0	0	1	0
individ	individual	0	0	1	1
säsongen	season	0	0	1	0
besluten	decisions	0	0	1	0
anus	ass	0	0	1	0
anus	anus	0	0	1	1
fysiska	natural	0	0	1	0
fysiska	physical	0	0	1	0
återstående	remaining	0	0	1	1
fysiskt	physically	0	0	1	1
fysiskt	physical	0	0	1	0
danny	danny	0	0	1	0
drevs	concentrated	0	0	1	0
drevs	was driven	0	0	1	0
beslutet	the decision	0	0	1	0
konkreta	specific	0	0	1	0
konkreta	concrete	0	0	1	0
fiender	enemies	0	0	1	0
fienden	enemy	0	0	1	0
fienden	the enemy	0	0	1	0
medlemmarna	members	0	0	1	0
medlemmarna	the members	0	0	1	0
lugn	calm	0	0	1	1
präglade	prague	0	0	1	0
präglade	the	0	0	1	0
präglade	characterized	0	0	1	0
ursäkt	excuse	0	0	1	1
ursäkt	apology	0	0	1	1
jordytan	earth's surface	0	0	1	0
jordytan	earth crust	0	0	1	0
fordon	vehicle/-s	0	0	1	0
fordon	vehicles	0	0	1	0
fordon	vehicle	0	0	1	1
genomförde	carried out	0	0	1	0
marklund	marklund	0	0	1	0
marijuana	marijuana	0	0	1	1
formerna	forms	0	0	1	0
träffades	met	0	0	1	0
träffades	was met	0	0	1	0
träffades	reached; met	0	0	1	0
regeringen	the government	0	0	1	0
regeringen	government	0	0	1	0
orsakerna	the causes	0	0	1	0
kevin	kevin	0	0	1	0
adeln	nobility	0	0	1	0
nikola	nikola	0	0	1	0
politiska	politic	0	0	1	0
politiska	political	0	0	1	0
påverkade	influenced	0	0	1	0
påverkade	affected	0	0	1	0
företeelse	experience; phenomenon; feature	0	0	1	0
företeelse	feature	0	0	1	0
företeelse	phenomenon	0	0	1	1
östtyskland	east germany	0	0	1	1
centralbanken	centralbank	0	0	1	0
centralbanken	central bank	0	0	1	0
potential	potential	0	0	1	0
politiskt	political	0	0	1	0
performance	performance	0	0	1	0
performance	uppträdande	0	0	1	0
centralstation	central station	0	0	1	0
magnetiska	magnetic	0	0	1	0
channel	channel	0	0	1	0
norman	norman	0	0	1	0
isolerad	isolation	0	0	1	0
isolerad	isolated	0	0	1	1
morden	murders	0	0	1	0
morden	the murders	0	0	1	0
förekommande	occuring	0	0	1	0
förekommande	where	0	0	1	0
fotografier	photographs	0	0	1	0
halvan	the half	0	0	1	0
halvan	half	0	0	1	0
politisk	political	0	0	1	1
beta	graze	0	0	1	1
beta	beta	0	0	1	1
mordet	the murder	0	0	1	0
mordet	murder	0	0	1	0
dahlén	dahlén	0	0	1	0
tränger	forces forward	0	0	1	0
tränger	cut in	0	0	1	0
tränger	penetration	0	0	1	0
japanerna	japanese	0	0	1	0
japanerna	the japanese	0	0	1	0
grundämne	elemental	0	0	1	0
grundämne	element	0	0	1	1
queens	queen	0	0	1	0
civilisationer	civilizations	0	0	1	0
otaliga	countless	0	0	1	0
otaliga	countless; endless	0	0	1	0
lojalitet	loyality	0	0	1	0
lojalitet	loyalty	0	0	1	1
påsk	easter	0	0	1	1
ämbetsmän	officers	0	0	1	0
ämbetsmän	bailies	0	0	1	0
ämbetsmän	officer	0	0	1	0
drottning	queen	0	0	1	1
allmänna	general	0	0	1	0
grammatik	grammar	0	0	1	1
framförde	performed	0	0	1	0
framförde	presented	0	0	1	0
kontrolleras	is controlled	0	0	1	0
kontrolleras	controlled	0	0	1	0
kontrollerar	controlling	0	0	1	0
kontrollerar	controls	0	0	1	0
kontrollerar	controls; controlling	0	0	1	0
ungdom	youth	0	0	1	1
civilisationen	civilization	0	0	1	0
härledas	derived	0	0	1	0
show	show	0	0	1	1
gränser	borders	0	0	1	0
gränser	frontiers	0	0	1	0
gränsen	border	0	0	1	0
gränsen	limit	0	0	1	0
gränsen	the line	0	0	1	0
adolfs	adolf's	0	0	1	0
adolfs	adolf	0	0	1	0
fånga	capture	0	0	1	1
fånga	capturing	0	0	1	0
tidigast	the earliest	0	0	1	0
führer	fuhrer	0	0	1	0
führer	fuehrer	0	0	1	0
generalsekreterare	the secretary-general	0	0	1	0
generalsekreterare	secretary general	0	0	1	1
samlingsalbum	compilation album	0	0	1	0
samlingsalbum	compilations	0	0	1	0
släktskap	relationship	0	0	1	1
släktskap	kinship	0	0	1	1
helig	holy	0	0	1	1
dick	dick	0	0	1	0
historier	stories	0	0	1	0
historier	history	0	0	1	0
jämförelse	comparative	0	0	1	0
jämförelse	comparison	0	0	1	1
jämförelse	jamfirelse	0	0	1	0
passande	fitting	0	0	1	1
passande	suitable	0	0	1	1
passande	matching	0	0	1	0
historien	history	0	0	1	1
diagnos	diagnostics	0	0	1	0
statsmakten	the government	0	0	1	0
statsmakten	power	0	0	1	0
statsmakten	government	0	0	1	0
förlorade	lost	0	0	1	0
karolinska	karolinska (institute for medicine)	0	0	1	0
karolinska	caroline	0	0	1	0
ges	given	0	0	1	0
ges	be given	0	0	1	0
ger	gives	0	0	1	0
ger	gives; is giving	0	0	1	0
ger	give	0	0	1	0
raser	races	0	0	1	0
raser	species	0	0	1	0
kulturellt	culture	0	0	1	0
kulturellt	cultural	0	0	1	0
kulturellt	culturally	0	0	1	0
konsolen	bracket	0	0	1	0
motsvarande	corresponding to	0	0	1	0
motsvarande	corresponding	0	0	1	1
källa	source	0	0	1	1
inspelningarna	recordings	0	0	1	0
kulturella	cultural	0	0	1	0
sällan	seldom	0	0	1	1
sällan	rare	0	0	1	0
katla	katla	0	0	1	0
katla	katla (fictive dragon in the classic "bröderna lejonhjärta")	0	0	1	0
vintergatan	milky way	0	0	1	1
vintergatan	the milky way	0	0	1	0
firade	celebrated	0	0	1	0
anklagelser	allegations	0	0	1	0
anklagelser	accusations	0	0	1	0
fortsättning	continuation	0	0	1	1
fortsättning	further accession	0	0	1	0
fortsättning	continued	0	0	1	0
gen	gene	0	0	1	1
beskyddare	protector	0	0	1	1
beskyddare	patron	0	0	1	1
himmlers	himmlers	0	0	1	0
himmlers	himmler	0	0	1	0
mattis	mattis	0	0	1	0
bengtsson	bengtsson	0	0	1	0
statistiska	statistical	0	0	1	0
förhindra	prevent	0	0	1	1
dianno	di'anno	0	0	1	0
dianno	dianno	0	0	1	0
spridda	spread	0	0	1	0
spridda	scattered	0	0	1	0
europacupen	euro (-pean) cup	0	0	1	0
europacupen	european cup	0	0	1	0
miley	miley	0	0	1	0
tolfte	twelth	0	0	1	0
tolfte	twelfth	0	0	1	1
relativt	relative	0	0	1	0
relativt	relatively	0	0	1	1
fokuserar	focuses	0	0	1	0
fokuserar	focus	0	0	1	0
nazisterna	the nazis	0	0	1	0
nazisterna	nazis	0	0	1	0
toppade	topped	0	0	1	0
teoretisk	theoretical	0	0	1	1
relativa	relative	0	0	1	0
sean	seab	0	0	1	0
sean	sean	0	0	1	0
stadsdelar	districts	0	0	1	0
stadsdelar	city districts	0	0	1	0
stadsdelar	neighborhoods	0	0	1	0
utgiven	published	0	0	1	0
menat	meant	0	0	1	0
menar	means	0	0	1	0
menar	mean	0	0	1	0
kandidater	candidates	0	0	1	0
stad	city	0	0	1	0
visades	was	0	0	1	0
visades	showed	0	0	1	0
vanns	was won	0	0	1	0
vanns	(was) won	0	0	1	0
bönor	beans	0	0	1	0
tränade	trained	0	0	1	0
bestämdes	was decided	0	0	1	0
bestämdes	decided	0	0	1	0
bestämdes	was determined	0	0	1	0
personligt	personal	0	0	1	0
personligt	private	0	0	1	0
gaga	gaga	0	0	1	0
personliga	personal	0	0	1	0
tsaren	the czar	0	0	1	0
tsaren	czar	0	0	1	0
tsaren	the tsar	0	0	1	0
august	august	0	0	1	0
ju	the	0	0	1	1
ju	the more	0	0	1	0
tur	turn	0	0	1	1
tur	tour	0	0	1	1
tur	luck	0	0	1	1
forskaren	researcher	0	0	1	0
jr	jr.	0	0	1	0
jr	junior	0	0	1	0
motsättningar	oppositions	0	0	1	0
motsättningar	contradictions	0	0	1	0
motsättningar	frictions; clashes	0	0	1	0
timme	hour	0	0	1	1
långfilm	feature film	0	0	1	0
långfilm	feature movie	0	0	1	0
tum	inch	0	0	1	1
tum	inches	0	0	1	0
signaler	signals	0	0	1	0
inbördes	relative	0	0	1	0
inbördes	intermutual	0	0	1	0
välgörenhet	charity	0	0	1	1
ja	yes	0	0	1	1
ministrar	ministers	0	0	1	0
tänder	teeth	0	0	1	0
rugby	american fotboll	0	0	1	0
rugby	rugby	0	0	1	1
utvalda	selected	0	0	1	0
utvalda	selected; chosen	0	0	1	0
medellivslängd	average lifespan	0	0	1	0
medellivslängd	life expectancy	0	0	1	0
tour	tour	0	0	1	0
paret	pair	0	0	1	0
paret	the couple	0	0	1	0
paret	parathyroid	0	0	1	0
följeslagare	companions	0	0	1	0
följeslagare	companion	0	0	1	1
naturresurser	natural resources	0	0	1	0
rösterna	votes	0	0	1	0
rösterna	the votes	0	0	1	0
tryck	press	0	0	1	0
tryck	pressure	0	0	1	1
tryck	print	0	0	1	1
vilja	will	0	0	1	1
vilja	like	0	0	1	0
cancer	cancer	0	0	1	1
statschefen	the head of state	0	0	1	0
statschefen	head of state	0	0	1	0
syntes	synthesis	0	0	1	1
ägnar	spend time	0	0	1	0
ägnar	dedicated	0	0	1	0
ägnar	spends time	0	0	1	0
grundare	founder	0	0	1	1
miljöproblem	environmental problem	0	0	1	0
miljöproblem	environmental problems	0	0	1	0
miljöproblem	enviormental problem	0	0	1	0
stängdes	closed	0	0	1	0
lexikon	lexicon	0	0	1	1
barry	barry	0	0	1	0
bildats	formed	0	0	1	0
bildats	had formed	0	0	1	0
bildats	created	0	0	1	0
kirsten	kirsten	0	0	1	0
kirsten	kristen	0	0	1	0
industrin	industry	0	0	1	0
utsatta	exposed	0	0	1	0
mars	march	0	0	1	1
måla	target	0	0	1	0
måla	grinding	0	0	1	0
marx	marx	0	0	1	0
mary	mary	0	0	1	0
kultur	culture	0	0	1	1
flaggan	the flag	0	0	1	0
flaggan	flag	0	0	1	0
cobain	cobain	0	0	1	0
partido	partido	0	0	1	0
avskaffa	abolish	0	0	1	1
bmi	bmi	0	0	1	0
spelfilmer	motion pictures	0	0	1	0
spelfilmer	feature film	0	0	1	0
spelfilmer	feature films	0	0	1	0
meningen	meningen	0	0	1	0
meningen	sense	0	0	1	0
påverkades	was affected by	0	0	1	0
påverkades	affected	0	0	1	0
fortsatt	further	0	0	1	1
fortsatt	continued	0	0	1	1
sound	sound	0	0	1	0
läs	read	0	0	1	0
läs	las	0	0	1	0
ständigt	always	0	0	1	1
ständigt	constant	0	0	1	0
trådlös	wireless	0	0	1	1
ständiga	permanent	0	0	1	0
ständiga	constant	0	0	1	0
dragit	drawn	0	0	1	0
dragit	dragged	0	0	1	0
dragit	preferred	0	0	1	0
uppstod	developed	0	0	1	0
uppstod	was	0	0	1	0
gånger	times	0	0	1	0
konstnär	artist	0	0	1	1
lät	made	0	0	1	0
lät	had	0	0	1	0
lät	sounded	0	0	1	0
sjöss	sea	0	0	1	0
övervikt	obesity	0	0	1	0
övervikt	overweight	0	0	1	1
nionde	ninth	0	0	1	1
sahara	sahara	0	0	1	0
uppmanade	urged	0	0	1	0
uppmanade	encouraged	0	0	1	0
liknande	similiar	0	0	1	0
liknande	similar	0	0	1	1
förband	units; formations; bound (themselves)	0	0	1	0
förband	bond	0	0	1	0
sydkorea	south koreans	0	0	1	0
sydkorea	south korea	0	0	1	1
gången	time	0	0	1	0
par	pair	0	0	1	1
upplagor	editions	0	0	1	0
upplagor	the edition	0	0	1	0
upplagor	issues	0	0	1	0
paz	paz	0	0	1	0
lava	lava	0	0	1	1
infödda	native	0	0	1	0
infödda	natives	0	0	1	1
pan	pan	0	0	1	0
samt	also	0	0	1	0
samt	as well as	0	0	1	0
tidvis	times	0	0	1	0
föreslagits	suggested	0	0	1	0
föreslagits	was suggested	0	0	1	0
föreslagits	been suggested	0	0	1	0
bistånd	aid	0	0	1	1
bistånd	assistance	0	0	1	1
säkerhetsråd	security	0	0	1	0
säkerhetsråd	security council	0	0	1	0
running	running	0	0	1	0
kuba	cubans	0	0	1	0
kuba	cuba	0	0	1	1
slåss	fight	0	0	1	1
teknisk	technical	0	0	1	1
markus	marcus	0	0	1	0
fattas	taken	0	0	1	0
bang	bang	0	0	1	0
wahlgren	wahlgren	0	0	1	0
välja	select	0	0	1	1
gates	gates	0	0	1	0
bebyggelse	settlements	0	0	1	0
bebyggelse	settlement	0	0	1	1
bebyggelse	habitation	0	0	1	1
privatliv	private	0	0	1	0
privatliv	privatitv	0	0	1	0
×	x	0	0	1	0
äkta	authentic	0	0	1	1
äkta	married	0	0	1	0
äkta	genuine	0	0	1	1
okända	unknown	0	0	1	0
säger	said	0	0	1	0
säger	says	0	0	1	0
säger	claims; says	0	0	1	0
säkert	securely	0	0	1	0
skapelse	creation	0	0	1	1
församlingen	parish	0	0	1	0
församlingen	congregation	0	0	1	0
byggnad	building	0	0	1	1
reaktioner	reactions	0	0	1	0
jakten	the hunt	0	0	1	0
jakten	hunt	0	0	1	0
ideologiskt	ideologically	0	0	1	0
ideologiskt	ideological	0	0	1	0
bowie	bowie	0	0	1	0
livstid	lifetime	0	0	1	1
livstid	life span	0	0	1	0
åter	again	0	0	1	1
åter	undertake	0	0	1	0
åter	ater	0	0	1	0
programledare	host	0	0	1	0
gotland	gotland	0	0	1	1
ideologiska	ideological	0	0	1	0
motverka	prevent	0	0	1	0
motverka	counteract	0	0	1	1
motverka	counter	0	0	1	0
erkänna	recognize	0	0	1	1
vintern	the winter	0	0	1	0
vintern	winter	0	0	1	0
schwarzenegger	schwarzenegger	0	0	1	0
underarten	subspecies	0	0	1	0
underarten	sub species	0	0	1	0
mor	mother	0	0	1	1
haft	had	0	0	1	0
behåller	retain	0	0	1	0
behåller	keeps	0	0	1	0
jakt	hunt	0	0	1	1
jakt	hunting	0	0	1	1
simmons	simmons	0	0	1	0
mon	mon	0	0	1	0
mångfald	diversity	0	0	1	1
mångfald	variety	0	0	1	0
underarter	sub-species	0	0	1	0
underarter	subspecies	0	0	1	0
baltiska	baltic	0	0	1	0
kollektiv	collective	0	0	1	1
kollektiv	public	0	0	1	0
mod	courage	0	0	1	1
mod	mod	0	0	1	0
christina	christina	0	0	1	0
adams	adams	0	0	1	0
manhattan	manhattan	0	0	1	0
km²	square kilometre	0	0	1	0
km²	kilometres	0	0	1	0
km²	km2	0	0	1	0
km²	km²	0	0	1	0
ställningar	positions	0	0	1	0
ställningar	standings	0	0	1	0
ställningar	notions	0	0	1	0
fångar	captures	0	0	1	0
fångar	prisoners	0	0	1	0
hög	high	0	0	1	1
hög	hog	0	0	1	0
rikskansler	chancellor	0	0	1	0
kategorisveriges	category sweden	0	0	1	0
hör	include	0	0	1	0
hör	belong	0	0	1	0
hör	hears	0	0	1	0
joan	joan	0	0	1	0
konspirationsteorier	conspiracy theories	0	0	1	0
jordbruket	agriculture	0	0	1	0
jordbruket	the agriculture	0	0	1	0
lotta	raffle	0	0	1	0
lotta	lotta	0	0	1	0
sudan	sudan	0	0	1	0
sudan	the sudan	0	0	1	0
löstes	solved	0	0	1	0
löstes	dissolved	0	0	1	0
drar	drag	0	0	1	0
drar	earn	0	0	1	0
övertygad	confident	0	0	1	0
övertygad	convinced	0	0	1	1
kmh	km/h	0	0	1	0
kmh	kmh	0	0	1	0
reportrar	reporters	0	0	1	0
konsten	art	0	0	1	0
konsten	the art	0	0	1	0
territorium	state	0	0	1	0
territorium	territory	0	0	1	1
samman	together	0	0	1	1
näringsliv	business	0	0	1	0
moderata	moderate	0	0	1	0
moderata	moderates	0	0	1	0
vistas	live	0	0	1	0
vistas	present	0	0	1	0
tunnlar	tunnels	0	0	1	0
londons	london's	0	0	1	0
cellen	cell	0	0	1	0
cellen	the cell	0	0	1	0
olof	olof	0	0	1	0
ifrågasatts	is questioned	0	0	1	0
ifrågasatts	questioned	0	0	1	0
ryggen	the back	0	0	1	0
ryggen	back	0	0	1	0
ändrades	changed	0	0	1	0
ändrades	was	0	0	1	0
tongivande	influential	0	0	1	0
marissa	marissa	0	0	1	0
tillverka	producing	0	0	1	0
celler	cells	0	0	1	0
östtysklands	east germany's	0	0	1	0
östtysklands	osttysklands	0	0	1	0
island	iceland	0	0	1	1
island	icelandic	0	0	1	0
förbjudet	prohibited	0	0	1	0
förbjuder	prohibiting	0	0	1	0
förbjuder	forbids	0	0	1	0
förbjuden	smoking	0	0	1	0
metaforer	metaphores	0	0	1	0
metaforer	metaphors	0	0	1	0
metaforer	metafor	0	0	1	0
lands	land	0	0	1	0
lands	on land	0	0	1	0
vanföreställningar	delusions	0	0	1	0
irländska	irish	0	0	1	0
lagarna	the laws	0	0	1	0
retoriken	rhetoric	0	0	1	0
auschwitz	auschwitz	0	0	1	0
sköta	manage	0	0	1	0
sköta	handle	0	0	1	0
sköta	operate	0	0	1	1
newtons	newton	0	0	1	0
newtons	newton's	0	0	1	0
wilde	wilde	0	0	1	0
beskrivas	described	0	0	1	0
beskrivas	be described	0	0	1	0
einstein	einstein	0	0	1	0
mark	soil	0	0	1	1
mark	territory	0	0	1	1
mark	ground	0	0	1	1
vindar	winds	0	0	1	0
fjädrar	spring	0	0	1	0
fjädrar	feathers	0	0	1	0
floderna	floods	0	0	1	0
floderna	the rivers	0	0	1	0
floderna	rivers	0	0	1	0
motivet	the motive	0	0	1	0
motivet	subject	0	0	1	0
behandling	treatment	0	0	1	1
varelse	creature	0	0	1	1
förhållande	in relation	0	0	1	0
förhållande	ratio	0	0	1	1
förhållande	(in) comparison (to)	0	0	1	0
anfalla	attack	0	0	1	1
uppskattades	estimated	0	0	1	0
uppskattades	appreciated	0	0	1	0
uppskattades	was appreciated	0	0	1	0
sålt	sold	0	0	1	0
omväxlande	varied	0	0	1	0
självt	itself	0	0	1	0
inletts	started	0	0	1	0
inletts	initiation	0	0	1	0
inletts	initiated	0	0	1	0
utbredd	widespread	0	0	1	1
utbredd	spread	0	0	1	1
själva	self	0	0	1	0
själva	actual	0	0	1	0
birger	birger	0	0	1	0
e	e	0	0	1	1
egen	own	0	0	1	1
arméns	the army's	0	0	1	0
arméns	arm	0	0	1	0
arméns	army's	0	0	1	0
woman	woman	0	0	1	0
mänsklig	human	0	0	1	1
världsturné	world tour	0	0	1	0
omröstning	vote	0	0	1	1
ronaldo	ronaldo	0	0	1	0
vhs	vhs	0	0	1	0
exemplar	copies	0	0	1	0
exemplar	example	0	0	1	1
bibliografi	bibliography	0	0	1	1
manuel	manuel	0	0	1	0
manuel	manual	0	0	1	0
verkliga	real	0	0	1	0
verkliga	fair	0	0	1	0
äta	eat	0	0	1	1
strömmar	flow	0	0	1	0
strömmar	streams	0	0	1	0
humanismen	humanism	0	0	1	0
parlament	parliament	0	0	1	1
youtube	youtube	0	0	1	0
manliga	male	0	0	1	0
populära	popular	0	0	1	0
deep	deep	0	0	1	0
general	general	0	0	1	1
skriven	written	0	0	1	1
pompejus	pompey	0	0	1	0
pompejus	pompejus	0	0	1	0
populärt	popular	0	0	1	0
populärt	popularly	0	0	1	1
erbjöd	offered	0	0	1	0
hästen	the horse	0	0	1	0
videon	the video	0	0	1	0
videon	video	0	0	1	0
film	film	0	0	1	1
again	again	0	0	1	0
genrer	genres	0	0	1	0
effekt	effect	0	0	1	1
effekt	power	0	0	1	1
istanbul	istanbul	0	0	1	1
rubiks	rubiks	0	0	1	0
rubiks	rubik's	0	0	1	0
muren	wall	0	0	1	0
förtryck	opression	0	0	1	0
kategorilevande	category of live	0	0	1	0
produktiv	productive	0	0	1	1
produktiv	productivity	0	0	1	0
stannade	stayed	0	0	1	0
behövde	did	0	0	1	0
behövde	needed	0	0	1	0
sammansättning	composition	0	0	1	1
genren	genre	0	0	1	0
faktorer	factors	0	0	1	0
rummet	room	0	0	1	0
ordna	arranging	0	0	1	0
ordna	arrange	0	0	1	1
profet	prophet	0	0	1	1
håkansson	hakansson	0	0	1	0
håkansson	håkansson	0	0	1	0
försvar	defence	0	0	1	1
försvar	defense	0	0	1	1
rykten	rumors	0	0	1	0
ledning	conduit	0	0	1	0
ledning	guidance	0	0	1	1
henriks	henry	0	0	1	0
kyros	cyrus	0	0	1	0
skapade	made	0	0	1	0
skapade	created	0	0	1	0
medicinska	medicinal	0	0	1	0
medicinska	medical	0	0	1	0
araberna	arabs	0	0	1	0
palestinska	palestinian	0	0	1	0
uppfostran	upbringing	0	0	1	1
u	u	0	0	1	0
dvs	(det vill säga) namely that	0	0	1	0
dvs	d.v.s.	0	0	1	0
dvs	i.e.	0	0	1	0
försörja	support	0	0	1	1
kuwait	kuwait	0	0	1	1
snabbaste	rapid	0	0	1	0
snabbaste	fastest	0	0	1	0
resolution	resolution	0	0	1	0
vila	rest	0	0	1	1
socialismen	the socialism	0	0	1	0
socialismen	socialism	0	0	1	0
inspirerat	inspired	0	0	1	0
dollar	dollar	0	0	1	1
vill	will	0	0	1	0
vill	to	0	0	1	0
vill	want	0	0	1	0
ström	power	0	0	1	0
ström	stream	0	0	1	1
ström	icon	0	0	1	0
hindrar	prevent	0	0	1	0
hindrar	stop; prevent	0	0	1	0
hindrar	prevents	0	0	1	0
skrivet	written	0	0	1	0
inspirerad	inspired	0	0	1	1
liam	liam	0	0	1	0
levern	the liver	0	0	1	0
levern	liver	0	0	1	0
sund	healthy	0	0	1	1
sund	narrow	0	0	1	0
sund	sane	0	0	1	1
världsliga	worldly	0	0	1	0
symbolen	the symbol	0	0	1	0
förbund	union	0	0	1	1
förbund	federal	0	0	1	0
förbund	league; alliance; union; compact; covenant	0	0	1	0
lugna	reassure	0	0	1	1
lugna	calm	0	0	1	1
indiska	indian	0	0	1	0
rwanda	rwanda	0	0	1	0
falska	fold	0	0	1	0
falska	false	0	0	1	0
symboler	symbols	0	0	1	0
skydda	protect	0	0	1	1
skydda	protection	0	0	1	0
skriver	write	0	0	1	0
skriver	type	0	0	1	0
seriens	series	0	0	1	0
kasta	discard	0	0	1	0
kasta	throw	0	0	1	1
utställning	display	0	0	1	1
utställning	exhibition	0	0	1	1
avhandling	treatise	0	0	1	1
avhandling	thesis	0	0	1	1
svår	severe	0	0	1	1
svår	difficult	0	0	1	1
handlade	dealt with	0	0	1	0
handlade	was (about); traded	0	0	1	0
handlade	was	0	0	1	0
israeliska	israeli	0	0	1	0
israeliska	isrealic	0	0	1	0
vägnät	network	0	0	1	0
ramen	frame	0	0	1	0
ramel	ramel	0	0	1	0
tät	compact	0	0	1	1
tät	frequent	0	0	1	1
tät	sealed	0	0	1	0
kulminerade	culminated	0	0	1	0
ansvarig	charge	0	0	1	0
långvariga	long-standing	0	0	1	0
långvariga	long	0	0	1	0
långvarigt	long-running	0	0	1	0
långvarigt	prolonged	0	0	1	0
långvarigt	long-standing	0	0	1	0
snuset	snuff	0	0	1	0
snuset	the snuff	0	0	1	0
säsonger	seasons	0	0	1	0
strålningen	the radiation	0	0	1	0
strålningen	radiation	0	0	1	0
suttit	been	0	0	1	0
suttit	sat	0	0	1	0
uppnår	reaches	0	0	1	0
uppnår	achieve	0	0	1	0
uppnås	obtained	0	0	1	0
uppnås	is achieved	0	0	1	0
ockuperades	occupied	0	0	1	0
cornelis	cornelis	0	0	1	0
lärare	teacher	0	0	1	1
sjönk	decreased	0	0	1	0
sjönk	sank	0	0	1	0
sjönk	sunk	0	0	1	0
massor	lots	0	0	1	0
massor	(in) masses	0	0	1	0
massor	tons	0	0	1	0
sjöng	sang	0	0	1	0
följde	followed	0	0	1	0
intressant	interestingly	0	0	1	1
intressant	of interest	0	0	1	0
håller	is	0	0	1	0
håller	holds	0	0	1	0
håller	halls	0	0	1	0
abc	abc (swedish news program)	0	0	1	0
abc	abc	0	0	1	1
hållet	attached via	0	0	1	0
hållet	cohesive	0	0	1	0
hållet	way	0	0	1	0
upphört	ceased	0	0	1	0
upphört	left the association	0	0	1	0
upphört	end	0	0	1	0
söder	south	0	0	1	1
danmark	denmark	0	0	1	1
uppståndelse	resurrection	0	0	1	1
publik	audience	0	0	1	1
publik	public	0	0	1	1
dvärghundar	miniature dogs	0	0	1	0
public	public	0	0	1	0
bebott	inhabit	0	0	1	0
bebott	inhabited	0	0	1	0
bebott	an inhabitated	0	0	1	0
vald	elected	0	0	1	0
vald	selected	0	0	1	1
jonas	jonas	0	0	1	0
kandidat	candidate	0	0	1	1
benen	legs	0	0	1	0
inställning	attitude	0	0	1	1
inställning	setting	0	0	1	0
inställning	view	0	0	1	0
fristående	independent	0	0	1	0
fristående	stand-alone	0	0	1	1
sistnämnda	later	0	0	1	0
sistnämnda	last	0	0	1	0
sistnämnda	sistamnda	0	0	1	0
vänta	(have to) wait; expect	0	0	1	0
vänta	wait	0	0	1	1
division	division	0	0	1	1
årsåldern	age group	0	0	1	0
årsåldern	years old	0	0	1	0
historiker	historians	0	0	1	0
jackie	jackie	0	0	1	0
airport	airport	0	0	1	0
förutsättningar	prerequisites	0	0	1	0
förutsättningar	(pre-)conditions	0	0	1	0
förutsättningar	condition	0	0	1	0
uppslagsverk	encyclopedia	0	0	1	0
uppslagsverk	encyklopedia	0	0	1	0
västerländska	vasterlandska	0	0	1	0
västerländska	western	0	0	1	0
amadeus	amadeus	0	0	1	0
alexandria	alexandria	0	0	1	0
utsträckning	extent	0	0	1	1
sjukhuset	the hospital	0	0	1	0
sjukhuset	hospital	0	0	1	0
africa	africa	0	0	1	0
förenklat	simplified	0	0	1	0
förenklat	made easier	0	0	1	0
enat	united	0	0	1	0
ocheller	and/or	0	0	1	0
hyllning	tribute	0	0	1	1
hyllning	tribute; homage	0	0	1	0
eye	eye	0	0	1	0
tävlade	competed	0	0	1	0
torrt	dry	0	0	1	0
besökte	visited	0	0	1	0
innebar	meant	0	0	1	0
innebar	was; meant; entailed	0	0	1	0
innebar	was	0	0	1	0
torra	dry	0	0	1	0
landet	state	0	0	1	0
landet	the country	0	0	1	0
diamond	diamond	0	0	1	0
leonard	leonard	0	0	1	0
koma	coma	0	0	1	1
brist	non	0	0	1	0
brist	lack	0	0	1	1
brist	failure; lack of	0	0	1	0
tillkommer	reside	0	0	1	0
tillkommer	will be	0	0	1	0
tillkommer	will be added	0	0	1	0
upptäckte	discovered	0	0	1	0
upptäckte	found	0	0	1	0
skivor	plates	0	0	1	0
skivor	records	0	0	1	0
förespråkar	occurring crackles	0	0	1	0
förespråkar	advocate	0	0	1	0
förespråkar	advocates	0	0	1	0
säker	items	0	0	1	0
säker	safe	0	0	1	1
säker	safety	0	0	1	0
vladimir	vladimir	0	0	1	0
tillverkningen	production	0	0	1	0
tillverkningen	the production	0	0	1	0
des	des	0	0	1	0
det	is	0	0	1	0
det	it	0	0	1	1
det	dent	0	0	1	0
roosevelt	roosevelt	0	0	1	0
del	part	0	0	1	1
lindgren	lindgren	0	0	1	0
den	it	0	0	1	1
befintliga	current	0	0	1	0
befintliga	existing	0	0	1	0
samtliga	all	0	0	1	1
hastigt	rapidly	0	0	1	1
hastigt	fast	0	0	1	1
förstaplatsen	first place	0	0	1	0
latinets	latin	0	0	1	0
latinets	the latin's	0	0	1	0
latinets	the latin	0	0	1	0
sovjetunionens	soviet union's; soviet's	0	0	1	0
sovjetunionens	soviet union	0	0	1	0
sugga	barrier	1	0	1	0
sugga	coins	1	0	1	0
sugga	soe	1	1	0	0
sugga	block	1	0	1	0
sugga	sow	1	1	0	1
betoning	stress	0	0	1	1
sjukdom	illness	0	0	1	1
sjukdom	disease	0	0	1	1
robinson	robinson	0	0	1	0
protein	protein	0	0	1	1
makten	power	0	0	1	0
makten	the power	0	0	1	0
stil	type	0	0	1	0
psykotiska	psychotic	0	0	1	0
varierat	varied	0	0	1	0
vänskap	friendship	0	0	1	1
stig	stig	0	0	1	0
stig	path	0	0	1	1
verkligheten	real	0	0	1	0
verkligheten	reality	0	0	1	0
dåliga	poor	0	0	1	0
dåliga	bad	0	0	1	0
blad	leaves	0	0	1	0
blad	leaf	0	0	1	1
undervisningen	teaching	0	0	1	0
undervisningen	the education	0	0	1	0
vikten	importance	0	0	1	0
vikten	weight	0	0	1	0
vikten	vikte	0	0	1	0
förekomst	presence	0	0	1	1
beteckna	denote the	0	0	1	0
beteckna	denote	0	0	1	1
makter	powers	0	0	1	0
sekulär	secular	0	0	1	1
rastafari	rastafari	0	0	1	0
rastafari	rastafarian	0	0	1	0
lina	line	0	0	1	1
lina	lina	0	0	1	0
engelske	the english	0	0	1	0
engelske	british	0	0	1	0
engelske	english	0	0	1	0
pettersson	pettersson	0	0	1	0
laboratorium	laboratory	0	0	1	1
judiska	jewish	0	0	1	0
motståndsrörelsen	the resistance	0	0	1	0
motståndsrörelsen	resistance	0	0	1	0
huvudkontor	central office	0	0	1	0
huvudkontor	headquarters	0	0	1	1
ligger	lies	0	0	1	0
ligger	is	0	0	1	0
påbörjas	start	0	0	1	0
påbörjas	begin	0	0	1	0
påbörjas	starts	0	0	1	0
vatten	water	0	0	1	1
rastafarianer	the rastafarian	0	0	1	0
rastafarianer	rastafarians	0	0	1	0
rastafarianer	rastafarian	0	0	1	0
rockgrupper	rock groups	0	0	1	0
rockgrupper	rock group	0	0	1	0
rockgrupper	rock bands	0	0	1	0
facebook	facebook	0	0	1	0
edwin	edwin	0	0	1	0
konservatismen	conservatism	0	0	1	0
civila	civil	0	0	1	0
bernadotte	bernadotte	0	0	1	0
uppgav	said	0	0	1	0
officiella	official	0	0	1	0
latinamerika	latin america	0	0	1	1
gradvis	gradually	0	0	1	1
gradvis	progressively	0	0	1	0
same	lapp	0	0	1	1
same	sami	0	0	1	0
sällsynta	rare	0	0	1	0
sydvästra	southwestern	0	0	1	0
sydvästra	southwest	0	0	1	0
diskussion	discussion	0	0	1	1
edmund	edmund	0	0	1	0
epok	epoch	0	0	1	1
gustafsson	gustafsson	0	0	1	0
saknades	lacked	0	0	1	0
saknades	missing	0	0	1	0
trossamfund	religious community	0	0	1	1
trossamfund	faith community	0	0	1	0
trossamfund	religious communities	0	0	1	0
områdena	the areas	0	0	1	0
områdena	areas	0	0	1	0
good	good	0	0	1	0
ängssyra	sorrel	1	1	0	1
ängssyra	suppress	1	0	1	0
ängssyra	Ängssyra	1	0	1	0
ängssyra	sorell	1	0	1	0
ängssyra	suppression	1	0	1	0
ängssyra	sorrels	1	0	1	0
ängssyra	angssyra (perennial herb)	1	0	1	0
egentliga	real one	0	0	1	0
egentliga	actual	0	0	1	0
fortsätta	remain	0	0	1	0
fortsätta	continue	0	0	1	1
oxford	oxford	0	0	1	1
skrifterna	scriptures	0	0	1	0
association	association	0	0	1	1
utöver	addition	0	0	1	0
porto	postage	0	0	1	1
robbie	bobbie	0	0	1	0
robbie	robbie	0	0	1	0
kungarna	the kings	0	0	1	0
kungarna	kings	0	0	1	0
namibia	namibia	0	0	1	0
tillträdde	assumed	0	0	1	0
tillträdde	took	0	0	1	0
tillträdde	tilltradde	0	0	1	0
out	out	0	0	1	0
inleder	start	0	0	1	0
inleder	initiates	0	0	1	0
haile	haile	0	0	1	0
genomgått	experienced	0	0	1	0
genomgått	passed	0	0	1	0
mental	mental	0	0	1	1
house	house	0	0	1	0
energy	energy	0	0	1	0
hard	hard	0	0	1	0
flytta	move	0	0	1	1
befäl	command	0	0	1	1
energi	energy	0	0	1	1
perry	perry	0	0	1	0
sanningen	truth	0	0	1	0
sanningen	the truth	0	0	1	0
förväntningar	expectations	0	0	1	0
oftast	usually	0	0	1	0
oftast	most often	0	0	1	0
infrastrukturen	infrastructure	0	0	1	0
infrastrukturen	the infrastructure	0	0	1	0
forskning	research	0	0	1	1
perro	perro	0	0	1	0
medför	means	0	0	1	0
medför	result	0	0	1	0
medför	entails	0	0	1	0
redan	already	0	0	1	1
redan	has already	0	0	1	0
däggdjuren	mammals	0	0	1	0
däggdjuren	the mammals	0	0	1	0
prins	prince	0	0	1	1
prins	prins	0	0	1	0
bönderna	the farmers	0	0	1	0
bönderna	farmers	0	0	1	0
lawrence	lawrence	0	0	1	0
eventuella	any	0	0	1	0
eventuella	eventual	0	0	1	0
blekinge	blekinge	0	0	1	0
uralbergen	the ural mountains	0	0	1	0
uralbergen	urals	0	0	1	0
uralbergen	ralbergen	0	0	1	0
eventuellt	possibly	0	0	1	1
eventuellt	eventually	0	0	1	0
viken	gulf	0	0	1	0
vägrade	refused	0	0	1	0
oklart	clear	0	0	1	0
inflationen	inflation	0	0	1	0
investeringar	investments	0	0	1	0
finland	finland	0	0	1	1
styrs	is controlled	0	0	1	0
styrs	ruled	0	0	1	0
tänkande	thinking	0	0	1	1
harris	harris	0	0	1	0
styre	rule	0	0	1	1
styre	governance	0	0	1	0
legenden	legend	0	0	1	0
ensam	alone	0	0	1	1
styra	controlling	0	0	1	0
styra	steer	0	0	1	1
top	top	0	0	1	0
färdig	pre	0	0	1	0
färdig	done	0	0	1	1
sjunkande	sinking; decreasing	0	0	1	0
sjunkande	decreasing	0	0	1	0
dont	do	0	0	1	0
saltkråkan	saltkrakan	0	0	1	0
saltkråkan	salt crow	0	0	1	0
något	any	0	0	1	1
något	something	0	0	1	1
råvaror	raw	0	0	1	0
råvaror	wood	0	0	1	0
råvaror	raw materials	0	0	1	0
snarast	rather	0	0	1	0
snarast	as soon as possible	0	0	1	0
carter	carter	0	0	1	0
kom	came	0	0	1	0
kol	charcoal	0	0	1	0
kol	coal; charcoal	0	0	1	0
kon	group	0	0	1	0
bay	bay	0	0	1	0
noga	carefully	0	0	1	0
observationer	observations	0	0	1	0
världens	the world's	0	0	1	0
världens	the world	0	0	1	0
världens	the worlds	0	0	1	0
möjlighet	an opportunity	0	0	1	0
möjlighet	oppertunity	0	0	1	0
möjlighet	possibility	0	0	1	1
kategoriasiens	category of asia	0	0	1	0
införts	been inserted	0	0	1	0
införts	introduced	0	0	1	0
kardinal	cardinal	0	0	1	1
samväldet	commonwealth	0	0	1	0
samväldet	the commonwealth	0	0	1	0
triangeln	triangle	0	0	1	0
triangeln	the triangle	0	0	1	0
part	party	0	0	1	1
gudarna	the gods	0	0	1	0
domstolen	court	0	0	1	0
domstolen	the court	0	0	1	0
matteusevangeliet	gospel of matthew	0	0	1	0
matteusevangeliet	book of matthew	0	0	1	0
också	also	0	0	1	1
fort	fast	0	0	1	1
fort	quickly	0	0	1	1
fattiga	poor	0	0	1	0
kväll	evening	0	0	1	1
upplysningen	the enlightenment	0	0	1	0
upplysningen	enlightenment	0	0	1	0
knapp	scarce	0	0	1	1
knapp	button	0	0	1	1
knapp	bare	0	0	1	0
proteinerna	the proteins	0	0	1	0
proteinerna	proteins	0	0	1	0
hämnd	revenge	0	0	1	1
nådde	reached	0	0	1	0
personens	person	0	0	1	0
personens	the persons	0	0	1	0
personens	the person's	0	0	1	0
älska	love	0	0	1	1
avtar	declines	0	0	1	0
avtar	avatar	0	0	1	0
avtar	decreases	0	0	1	0
lyssnar	listens	0	0	1	0
lyssnar	listen	0	0	1	0
rikedom	riches	0	0	1	1
rikedom	wealth	0	0	1	1
militärt	military	0	0	1	0
militärt	militarily	0	0	1	0
årtionde	decade	0	0	1	1
gjord	made	0	0	1	1
militära	military	0	0	1	0
någon	someone	0	0	1	1
någon	anybody	0	0	1	1
rättegång	trial	0	0	1	1
rättegång	steering wheel gang	0	0	1	0
flertalet	most	0	0	1	0
flertalet	several	0	0	1	0
flertalet	majority; plurality	0	0	1	0
gjort	made	0	0	1	0
gjort	done	0	0	1	1
gjort	created	0	0	1	0
mountain	mountain	0	0	1	0
hundratals	hundreds of	0	0	1	0
hundratals	hundreds	0	0	1	0
svagare	weaker	0	0	1	0
svagare	weak	0	0	1	0
sång	song	0	0	1	1
gärdestad	nugent	0	0	1	0
gärdestad	garden city	0	0	1	0
caesar	caesar	0	0	1	0
genast	at once	0	0	1	1
genast	immediately	0	0	1	1
taktik	tactics	0	0	1	1
taktik	tactic	0	0	1	0
taktik	strategy	0	0	1	0
inkomsterna	the incomes	0	0	1	0
inkomsterna	the income	0	0	1	0
inkomsterna	revenue	0	0	1	0
skjuta	delay	0	0	1	0
skjuta	postpone; shoot	0	0	1	0
patterson	patterson	0	0	1	0
krafter	forces	0	0	1	0
gillade	liked	0	0	1	0
gillade	approved; liked	0	0	1	0
niclas	niclas	0	0	1	0
kraften	the force	0	0	1	0
kraften	power	0	0	1	0
identifiera	identification	0	0	1	0
utbrott	outbreak	0	0	1	1
utbrott	outbreaks	0	0	1	0
samtidigt	while	0	0	1	0
samtidigt	simultaneous	0	0	1	0
organiserade	organized	0	0	1	0
kända	known	0	0	1	0
tvärtom	on the contrary	0	0	1	1
tvärtom	contrary to	0	0	1	0
tvärtom	vice versa	0	0	1	0
ko	co	0	0	1	0
ko	cow	0	0	1	1
varför	therefore	0	0	1	0
varför	why did	0	0	1	0
varför	why	0	0	1	1
km	km	0	0	1	0
km	kilometers	0	0	1	0
kl	hr	0	0	1	0
kl	at	0	0	1	0
kl	o'clock	0	0	1	0
kr	kronas	0	0	1	0
liechtenstein	liechtenstein	0	0	1	0
hända	may	0	0	1	0
hända	provide	0	0	1	0
organism	organism	0	0	1	1
hände	happened	0	0	1	1
thomas	thomas	0	0	1	0
venedig	venice	0	0	1	0
venedig	venedig	0	0	1	0
kvalitet	kvalilet	0	0	1	0
kvalitet	quality	0	0	1	1
tillhör	belongs	0	0	1	0
tillhör	belonging to	0	0	1	0
byttes	changed	0	0	1	0
byttes	was exchanged	0	0	1	0
relation	ratio	0	0	1	0
relation	relation	0	0	1	1
utveckla	develop	0	0	1	1
utveckla	developing	0	0	1	0
fina	beautiful	0	0	1	0
fina	fine	0	0	1	0
valet	selection	0	0	1	0
valet	the election	0	0	1	0
antagit	adopted	0	0	1	0
antagit	presumed	0	0	1	0
hänsyn	light	0	0	1	0
hänsyn	consideration	0	0	1	1
kristna	christian	0	0	1	0
reaktionen	reaction	0	0	1	0
reaktionen	the reaction	0	0	1	0
plötsligt	suddenly	0	0	1	1
plötsligt	sudden	0	0	1	0
wallenberg	wallenberg	0	0	1	0
röd	rod	0	0	1	0
röd	red	0	0	1	1
medverka	take part	0	0	1	1
medverka	participate	0	0	1	0
tionde	tenth	0	0	1	1
karaktäriseras	characterizes	0	0	1	0
karaktäriseras	is characterised	0	0	1	0
karaktäriseras	is charactarized	0	0	1	0
avseende	regard	0	0	1	1
avseende	for	0	0	1	0
förena	combine	0	0	1	1
förena	unite	0	0	1	1
förena	combining	0	0	1	0
blomstrade	flourished	0	0	1	0
fröväxter	about	1	0	1	0
fröväxter	seed-bearing plants	1	1	0	0
fröväxter	provaxter	1	0	1	0
fröväxter	seed plants	1	1	0	0
fröväxter	phanerogams	1	0	1	0
fröväxter	seed plant	1	1	0	0
fröväxter	seedlings	1	0	1	0
fröväxter	spermatophytes	1	0	1	0
fröväxter	spermatophyte	1	1	0	0
fröväxter	with	1	0	1	0
notation	notation	0	0	1	0
beslutar	decides	0	0	1	0
express	express	0	0	1	1
beslutat	resolved	0	0	1	0
beslutat	decided	0	0	1	0
typiska	typical	0	0	1	0
husen	housing	0	0	1	0
husen	the houses	0	0	1	0
erkännande	recognition	0	0	1	0
sänker	lowers	0	0	1	0
sänker	lower	0	0	1	0
sänker	sinks	0	0	1	0
rör	touch	0	0	1	0
rör	touches	0	0	1	0
rör	move(-s)	0	0	1	0
rör	row	0	0	1	0
wallander	wallander	0	0	1	0
gamle	old	0	0	1	0
tjänster	services	0	0	1	0
uttrycket	the expression	0	0	1	0
uttrycket	expression	0	0	1	0
uttrycker	express	0	0	1	0
uttrycker	expressing	0	0	1	0
uttrycker	express (-es)	0	0	1	0
flykt	flight	0	0	1	1
flykt	escape	0	0	1	1
huset	housing	0	0	1	0
huset	the house	0	0	1	0
svarar	responds	0	0	1	0
somrar	summers	0	0	1	0
stadium	stage	0	0	1	0
styrdes	was guided	0	0	1	0
styrdes	governed	0	0	1	0
styrdes	ruled	0	0	1	0
tillhöra	belong to	0	0	1	1
tillhöra	belonging to	0	0	1	0
röst	voice	0	0	1	1
rollfigur	character	0	0	1	0
två	two	0	0	1	1
tengil	tengil	0	0	1	0
tillhört	belonged	0	0	1	0
tillhört	belonged to	0	0	1	0
båten	vessel	0	0	1	0
båten	the boat	0	0	1	0
båten	boat	0	0	1	0
rovdjur	predator	0	0	1	1
rovdjur	predators	0	0	1	0
fans	fans	0	0	1	0
upphör	end	0	0	1	0
landsbygden	rural	0	0	1	0
landsbygden	rural area	0	0	1	0
champagne	champagne	0	0	1	1
liberaler	liberals	0	0	1	0
romarriket	roman empire	0	0	1	0
romarriket	the roman empire	0	0	1	0
bildandet	setting-up	0	0	1	0
bildandet	establishment	0	0	1	0
bildandet	formation	0	0	1	0
professionella	professional	0	0	1	0
förklarades	was explained	0	0	1	0
förklarades	explained	0	0	1	0
kritiserades	critisized	0	0	1	0
kritiserades	critizised	0	0	1	0
skivorna	the records	0	0	1	0
skivorna	records	0	0	1	0
skivorna	plates	0	0	1	0
marilyn	marilyn	0	0	1	0
framställning	preparation	0	0	1	0
framställning	production	0	0	1	1
musklerna	muscles	0	0	1	0
musklerna	the muscles	0	0	1	0
statligt	state	0	0	1	0
statligt	governmental	0	0	1	0
erbjöds	offered	0	0	1	0
akon	akon	0	0	1	0
vuxit	grown	0	0	1	0
statliga	state	0	0	1	0
restaurang	restaurang	0	0	1	0
restaurang	restaurant	0	0	1	1
framförts	forward	0	0	1	0
framförts	performed	0	0	1	0
baltimore	baltimore	0	0	1	0
romska	romani	0	0	1	0
romska	roma	0	0	1	0
globala	global	0	0	1	0
kroatiens	croatia's	0	0	1	0
kroatiens	croatias	0	0	1	0
kroatiens	croatian	0	0	1	0
point	point	0	0	1	0
folkmord	genocide	0	0	1	1
andas	breath	0	0	1	1
andas	breathes	0	0	1	0
tennessee	tennessee	0	0	1	0
globalt	globally	0	0	1	0
globalt	global	0	0	1	0
inrättades	established	0	0	1	0
inrättades	were implemented	0	0	1	0
västergötland	västergötland	0	0	1	0
lyfta	lift	0	0	1	1
övertog	took over	0	0	1	0
övertog	overtook	0	0	1	0
laos	laos	0	0	1	0
förföljelser	persecution	0	0	1	0
förföljelser	pursuits	0	0	1	0
förföljelser	persecutions	0	0	1	0
förhandlingarna	the negotiations	0	0	1	0
förhandlingarna	negotiations	0	0	1	0
bengt	bengt	0	0	1	0
popularitet	popularity	0	0	1	1
gav	gave	0	0	1	0
effektiva	effective	0	0	1	0
gas	gas	0	0	1	1
besöka	visit	0	0	1	1
vana	familiar	0	0	1	0
vana	used	0	0	1	0
vana	habit	0	0	1	1
kalmar	kalmar	0	0	1	0
besökt	visited	0	0	1	0
effektivt	effective	0	0	1	0
trupperna	troops	0	0	1	0
trupperna	the troops	0	0	1	0
detsamma	the same	0	0	1	1
detsamma	same	0	0	1	0
bild	picture	0	0	1	1
bild	image	0	0	1	1
spridning	diffusion	0	0	1	1
spridning	distribution	0	0	1	1
spridning	proliferation	0	0	1	1
bill	car	0	0	1	0
villkoren	the terms	0	0	1	0
villkoren	conditions	0	0	1	0
religiösa	religious	0	0	1	0
portugal	portugal	0	0	1	1
arenan	arena	0	0	1	0
arenan	the arena	0	0	1	0
elektronik	electronics	0	0	1	1
släppas	released	0	0	1	0
släppas	be released	0	0	1	0
övers	transl	0	0	1	0
övers	translation	0	0	1	0
monroe	monroe - it's a persons name	0	0	1	0
monroe	monroe	0	0	1	0
rederiet	the shipping company	0	0	1	0
rederiet	the company	0	0	1	0
rederiet	shipping company	0	0	1	0
granska	examining	0	0	1	0
granska	review	0	0	1	1
granska	exam	0	0	1	0
sjuk	ill	0	0	1	1
sjuk	disease	0	0	1	0
hamna	end up	0	0	1	0
hamna	end	0	0	1	0
belägg	coating	0	0	1	0
belägg	evidence	0	0	1	1
administrationen	administration	0	0	1	0
förklara	explain	0	0	1	1
förklara	declaring	0	0	1	0
sittande	fitting	0	0	1	0
sittande	appointed	0	0	1	0
sittande	sitting	0	0	1	1
development	development	0	0	1	0
utmed	along	0	0	1	1
avrättade	executed	0	0	1	0
skotska	scotland	0	0	1	0
skotska	scottish	0	0	1	0
syd	south	0	0	1	1
fågelarter	bird species	0	0	1	0
fågelarter	species of bird	0	0	1	0
syn	sight	0	0	1	1
syn	view	0	0	1	1
jerusalems	jerusalem's	0	0	1	0
moment	step	0	0	1	0
kallades	was called	0	0	1	0
kallades	called	0	0	1	0
kallades	summoned	0	0	1	0
parentes	brackets	0	0	1	0
undersökningar	surveys; investigations	0	0	1	0
undersökningar	studies	0	0	1	0
undersökningar	studies'	0	0	1	0
mot	against	0	0	1	1
kungariket	kingdom	0	0	1	0
kungariket	the kingdom	0	0	1	0
engelsmännen	the british	0	0	1	0
engelsmännen	the english	0	0	1	0
engelsmännen	english people	0	0	1	0
noll	zero	0	0	1	1
kapitel	chapter	0	0	1	1
albanien	albania	0	0	1	1
jorderosion	earth erosion	0	0	1	0
jorderosion	soil erosion	0	0	1	0
åttonde	eighth	0	0	1	1
åttonde	the eighth	0	0	1	0
förståelse	understanding	0	0	1	1
colorblack	color black	0	0	1	0
skott	bulkheads	0	0	1	0
skott	round	0	0	1	0
skott	shots	0	0	1	0
albanska	albanian	0	0	1	0
norrland	northern	0	0	1	0
norrland	norrland	0	0	1	0
gränsar	border	0	0	1	0
gränsar	adjacent	0	0	1	0
gränsar	borders (to)	0	0	1	0
dikter	poems	0	0	1	0
bibeln	bible	0	0	1	0
kommunister	communists	0	0	1	0
juventus	juventus	0	0	1	0
halvt	half	0	0	1	1
organization	organization	0	0	1	0
representanter	represenatives	0	0	1	0
representanter	representatives	0	0	1	0
passerar	passes	0	0	1	0
passerar	pass	0	0	1	0
struktur	structure	0	0	1	1
senaste	last	0	0	1	0
alternativt	alternatively	0	0	1	0
alternativt	alternative	0	0	1	0
självständigheten	independance	0	0	1	0
självständigheten	independence	0	0	1	0
östtimor	east timor	0	0	1	0
world	world	0	0	1	0
hennes	her	0	0	1	1
analytiska	analytical	0	0	1	0
alternativa	alternative	0	0	1	0
förhandla	negotiate	0	0	1	1
förhandla	negotiating	0	0	1	0
sektion	section	0	0	1	1
tänkare	thinker	0	0	1	1
sparta	spartans	0	0	1	0
sparta	sparta	0	0	1	0
administrativt	administrative	0	0	1	0
administrativt	administratively	0	0	1	0
monarkin	monarchy	0	0	1	0
monarkin	the monarchy	0	0	1	0
administrativa	administrative	0	0	1	0
administrativa	administration	0	0	1	0
administrativa	administative	0	0	1	0
högste	supreme	0	0	1	0
högste	highest	0	0	1	0
högste	chief	0	0	1	0
högsta	highest	0	0	1	1
bin	bin	0	0	1	0
dubbelt	double	0	0	1	1
bil	car	0	0	1	1
teknik	technique	0	0	1	1
teknik	technology	0	0	1	0
teknik	technic	0	0	1	0
big	big	0	0	1	0
kejsaren	emperor	0	0	1	0
kejsaren	the emperor	0	0	1	0
avlidna	diseased	0	0	1	0
avlidna	deceased	0	0	1	0
avlidna	the perished	0	0	1	0
af	of	0	0	1	0
af	of (old swedish)	0	0	1	0
företeelser	phenomena	0	0	1	0
bit	piece	0	0	1	1
indonesiska	indonesian	0	0	1	0
utöva	carry	0	0	1	0
utöva	utÖva	0	0	1	0
utöva	exercise	0	0	1	1
kolonialtiden	the colonial times	0	0	1	0
kolonialtiden	colonial period	0	0	1	0
emigrerade	emigrated	0	0	1	0
terräng	off	0	0	1	0
terräng	terrain	0	0	1	1
människorna	men	0	0	1	0
människorna	the humans	0	0	1	0
princip	principle	0	0	1	1
princip	principal	0	0	1	0
använt	using	0	0	1	0
använt	used	0	0	1	0
vägg	wall	0	0	1	1
försökte	try	0	0	1	0
försökte	tried to	0	0	1	0
försökte	tried	0	0	1	1
anatomi	anatomy	0	0	1	1
google	google	0	0	1	0
stött	met	0	0	1	0
stött	supported	0	0	1	0
stött	stott	0	0	1	0
identisk	identical	0	0	1	1
egyptiska	egyptian	0	0	1	0
tolkningar	interpretations	0	0	1	0
tolkningar	interpretation	0	0	1	0
back	reverse	0	0	1	1
historisk	historic	0	0	1	1
historisk	historical	0	0	1	1
cocacola	coca cola	0	0	1	0
cocacola	coca-cola	0	0	1	0
lars	lars	0	0	1	0
flygplatser	airports	0	0	1	0
flygplatser	air ports	0	0	1	0
berättelsen	story	0	0	1	0
berättelsen	the story	0	0	1	0
integration	integration	0	0	1	1
per	per	0	0	1	1
pratar	talks	0	0	1	0
pratar	talking	0	0	1	0
pratar	talk	0	0	1	0
diplomatiska	diplomatic	0	0	1	0
saab	saab	0	0	1	0
enklare	easier	0	0	1	0
enklare	simpler	0	0	1	0
utgöra	compose	0	0	1	1
utgöra	make up	0	0	1	1
nordamerika	north america	0	0	1	1
överlevande	survivors	0	0	1	0
överlevande	over living	0	0	1	0
överlevande	survivor; survivors; surviving	0	0	1	0
vänstra	left-hand	0	0	1	0
vänstra	left	0	0	1	0
vasaloppet	vasaloppet	0	0	1	0
välkänd	known	0	0	1	0
välkänd	well-known	0	0	1	1
välkänd	well known	0	0	1	0
ockuperade	occupied	0	0	1	1
nödvändigt	neccessary	0	0	1	0
nödvändigt	necessary	0	0	1	0
britannica	britannica	0	0	1	0
korta	short	0	0	1	0
avlägsna	distant	0	0	1	0
avlägsna	remove	0	0	1	1
nödvändiga	necessary	0	0	1	0
nödvändiga	essential	0	0	1	0
fallit	fallen	0	0	1	0
fallit	fall	0	0	1	0
jimmy	jimmy	0	0	1	0
grammy	grammy	0	0	1	0
styrelse	government; direction	0	0	1	0
styrelse	board	0	0	1	1
styrelse	board of directors	0	0	1	0
barcelonas	barcelona	0	0	1	0
barcelonas	barcelona's	0	0	1	0
jobbar	work	0	0	1	0
jobbar	does the work	0	0	1	0
steven	steven	0	0	1	0
våren	spring	0	0	1	0
våren	the spring	0	0	1	0
ordnar	fix	0	0	1	0
ordnar	decorations	0	0	1	0
ordnar	arrange	0	0	1	0
författarskap	the writer	0	0	1	0
författarskap	authorship	0	0	1	1
ontario	ontario	0	0	1	0
förödande	devastating	0	0	1	1
ansvar	responsibilities	0	0	1	0
ansvar	responsibility	0	0	1	1
förre	pre	0	0	1	0
förre	former	0	0	1	1
förre	forrester	0	0	1	0
motståndarna	the opponents	0	0	1	0
motståndarna	opponents	0	0	1	0
förra	last	0	0	1	1
förra	former	0	0	1	1
turkiska	turkey	0	0	1	0
turkiska	turkish	0	0	1	1
berömda	famous	0	0	1	0
berömda	forceps	0	0	1	0
medvetande	awareness	0	0	1	0
medvetande	consciousnesses extensive	0	0	1	0
medvetande	consciousness	0	0	1	1
jaga	course	0	0	1	1
jaga	hunt	0	0	1	1
jaga	chase	0	0	1	1
serie	comic; row; succession; serial	0	0	1	0
serie	cartoon	0	0	1	0
serie	series	0	0	1	1
konsul	consulting	0	0	1	0
konsul	consul	0	0	1	1
utlösning	release	0	0	1	1
utlösning	ejaculation	0	0	1	0
utlösning	trigger	0	0	1	0
motståndare	opponent	0	0	1	1
motståndare	opponents	0	0	1	1
köpmän	traders	0	0	1	0
köpmän	merchants	0	0	1	0
torsten	torsten	0	0	1	0
jonathan	jonathan	0	0	1	0
skillnaden	the difference	0	0	1	0
göteborgs	gothenburgs	0	0	1	0
göteborgs	gothenburg	0	0	1	0
ledningen	conduit	0	0	1	0
ledningen	the lead	0	0	1	0
planen	the field	0	0	1	0
planen	the plan	0	0	1	0
planen	plan	0	0	1	0
planet	planet	0	0	1	1
smycken	jewlery	0	0	1	0
smycken	jewellery	0	0	1	0
litterär	literary	0	0	1	1
sultanen	sultan	0	0	1	0
planer	plans	0	0	1	0
amfetamin	amphetamine	0	0	1	1
skillnader	differences	0	0	1	0
reggaen	reggae	0	0	1	0
reggaen	the reggae	0	0	1	0
ställningen	position	0	0	1	0
reidar	reidar	0	0	1	0
titel	title	0	0	1	1
expedition	caretaker	0	0	1	0
expedition	expidition	0	0	1	0
expedition	expedition	0	0	1	1
kommittén	the committee	0	0	1	0
kommittén	committee	0	0	1	0
tropiskt	tropical	0	0	1	0
utförda	formed	0	0	1	0
utförda	performed	0	0	1	0
utförda	made	0	0	1	0
tropiska	tropical	0	0	1	0
tropiska	tropic	0	0	1	0
överföras	transfer	0	0	1	0
överföras	transferred	0	0	1	0
utförde	did	0	0	1	0
materia	matter	0	0	1	1
materia	materia	0	0	1	0
tyskland	germany	0	0	1	1
eller	or	0	0	1	1
voltaire	voltaire	0	0	1	0
familjer	families	0	0	1	0
familjen	the family	0	0	1	0
familjen	family	0	0	1	0
betalar	paying	0	0	1	0
betalar	pay	0	0	1	0
makedonien	macedonia	0	0	1	0
oerhörd	tremendous	0	0	1	0
anser	view	0	0	1	0
anser	believes	0	0	1	0
anses	be	0	0	1	0
anses	deemed; regarded	0	0	1	0
inåt	inwards	0	0	1	1
inåt	inwardly	0	0	1	0
ovanpå	top	0	0	1	0
ovanpå	on top of	0	0	1	0
maos	maos	0	0	1	0
maos	mao	0	0	1	0
maos	mao's	0	0	1	0
lena	lena	0	0	1	0
utvecklade	developed	0	0	1	0
utvecklade	oral	0	0	1	0
sekulära	secular	0	0	1	0
samla	collecting	0	0	1	0
samla	collect	0	0	1	1
samla	gather	0	0	1	1
mutationer	mutations	0	0	1	0
miljön	environment	0	0	1	0
miljön	the environment	0	0	1	0
skådespelare	actor	0	0	1	1
skådespelare	period players	0	0	1	0
nedgång	decline	0	0	1	1
nedgång	decreases	0	0	1	0
nedgång	fall	0	0	1	1
ritualer	rituals	0	0	1	0
storkors	the grand cross	0	0	1	0
talades	spoken	0	0	1	0
talades	spoken (of)	0	0	1	0
talades	spoke	0	0	1	0
regionala	regional	0	0	1	0
sambandet	the connection	0	0	1	0
sambandet	connection	0	0	1	0
sambandet	relation	0	0	1	0
dramatiker	playwright	0	0	1	0
dramatiker	dramatist	0	0	1	1
dramatiker	dramatists	0	0	1	0
judisk	jewish	0	0	1	1
judisk	jew	0	0	1	1
hertig	duke	0	0	1	1
regionalt	regional	0	0	1	0
regionalt	regionally	0	0	1	0
födelse	date	0	0	1	0
födelse	birth	0	0	1	1
flod	basin	0	0	1	0
flod	river	0	0	1	1
jason	jason	0	0	1	0
ökning	increase	0	0	1	1
tillgångar	assets	0	0	1	1
östblocket	east block	0	0	1	0
östblocket	the eastern bloc	0	0	1	0
östblocket	cheese block	0	0	1	0
stred	fought	0	0	1	0
uran	uranium	0	0	1	1
frankrike	france	0	0	1	1
dyrare	more expensive	0	0	1	0
dyrare	expensive	0	0	1	0
präster	priests	0	0	1	0
sigmund	sigmund	0	0	1	0
intensivt	intensive	0	0	1	0
intensivt	hard	0	0	1	0
privat	private	0	0	1	1
lilla	small	0	0	1	1
hindra	hinder	0	0	1	1
hindra	prevent	0	0	1	0
hindra	stop	0	0	1	0
medlemskap	membership	0	0	1	1
betrakta	view; regard	0	0	1	0
betrakta	view	0	0	1	1
sydafrikanska	south african	0	0	1	0
sydafrikanska	african	0	0	1	0
sahlin	sahlin	0	0	1	0
intensiva	intensive	0	0	1	0
intensiva	intense	0	0	1	0
kärnan	core	0	0	1	0
kärnan	the core	0	0	1	0
kollaps	collapse	0	0	1	1
atlas	atlas	0	0	1	1
graven	the grave	0	0	1	0
graven	grave	0	0	1	0
passiv	passive	0	0	1	1
huvudstaden	capital	0	0	1	0
kampanjen	campaign	0	0	1	0
plikt	duty	0	0	1	1
avgörande	settling	0	0	1	0
avgörande	decisive	0	0	1	1
avgörande	essential	0	0	1	0
stål	steel	0	0	1	1
stål	rate	0	0	1	0
annika	annika	0	0	1	0
varnade	warned	0	0	1	0
öns	the islands	0	0	1	0
öns	island's	0	0	1	0
utgjordes	was	0	0	1	0
utgjordes	make up	0	0	1	0
utgjordes	comprised; consisted	0	0	1	0
svts	svt	0	0	1	0
svts	svts	0	0	1	0
rede	coated	1	0	1	0
rede	network	1	1	0	0
rede	ways	1	0	1	0
rede	clutch	1	0	1	0
rede	nest	1	1	0	1
rede	means of	1	0	1	0
demokratisk	democratic	0	0	1	1
exemplet	the example	0	0	1	0
exemplet	example	0	0	1	0
säte	sate	0	0	1	0
säte	seat	0	0	1	1
knight	knight	0	0	1	1
joel	joel	0	0	1	0
dinosaurierna	dinosaurs	0	0	1	0
dinosaurierna	dinasaurs	0	0	1	0
sätt	manner	0	0	1	1
sätt	way	0	0	1	1
warszawa	warzaw	0	0	1	0
warszawa	warsaw	0	0	1	1
naturens	nature	0	0	1	0
naturens	nature's	0	0	1	0
joey	joey	0	0	1	0
fördragen	treaties	0	0	1	0
fördragen	the compacts	0	0	1	0
litterära	literary	0	0	1	0
litterära	literal	0	0	1	0
utbredda	widespread	0	0	1	0
utbredda	spread	0	0	1	0
vanligaste	frequent	0	0	1	0
vanligaste	most common	0	0	1	0
irländsk	irish	0	0	1	1
irländsk	ireland	0	0	1	0
strömning	strom accession	0	0	1	0
strömning	flow	0	0	1	0
carlo	carlo	0	0	1	0
depression	depression	0	0	1	1
fortsättningen	the continuation	0	0	1	0
fortsättningen	remain	0	0	1	0
övertala	convince	0	0	1	0
övertala	persuade	0	0	1	1
edison	edison	0	0	1	0
litteraturen	literature	0	0	1	0
mozarts	mozart	0	0	1	0
mozarts	mozart's	0	0	1	0
tillkomst	origin	0	0	1	1
tillkomst	established	0	0	1	0
tillkomst	advent	0	0	1	0
öppnade	opened	0	0	1	0
öppnade	opening	0	0	1	0
senare	latterly; later	0	0	1	0
senare	later	0	0	1	1
placering	position	0	0	1	0
placering	placement	0	0	1	0
analsex	analsex	0	0	1	0
analsex	anal sex	0	0	1	0
och	and	0	0	1	1
kyrka	church	0	0	1	1
extremt	extremely	0	0	1	0
extremt	extreme angular	0	0	1	0
extremt	extreme	0	0	1	0
luis	luis	0	0	1	0
extrema	extreme	0	0	1	0
sina	their	0	0	1	0
sina	his	0	0	1	0
honom	his	0	0	1	0
honom	him	0	0	1	1
medeltid	medieval	0	0	1	0
medeltid	the medieval times	0	0	1	0
arbetslöshet	unemplyment	0	0	1	0
arbetslöshet	unemployment	0	0	1	1
turkar	turks	0	0	1	0
alaska	alaska	0	0	1	1
sällsynt	rare	0	0	1	1
omgången	round	0	0	1	0
lagts	added	0	0	1	0
katolicismen	catholisism	0	0	1	0
katolicismen	catholicism	0	0	1	0
underhåll	support	0	0	1	1
underhåll	allowance	0	0	1	1
underhåll	entertainment	0	0	1	0
miljard	billion	0	0	1	1
miljard	one billion	0	0	1	0
uranus	uranus	0	0	1	1
honor	ära	0	0	1	0
honor	female	0	0	1	0
existens	existence	0	0	1	1
protokoll	protocol	0	0	1	1
talare	speakers	0	0	1	0
talare	speaker	0	0	1	1
talare	spoke	0	0	1	0
privata	private	0	0	1	0
stundom	sometimes	0	0	1	1
stundom	somtimes	0	0	1	0
filippinerna	filipinos	0	0	1	0
filippinerna	the philippines	0	0	1	0
betraktas	considered	0	0	1	0
betraktar	regard	0	0	1	0
betraktar	sees	0	0	1	0
ovan	above	0	0	1	1
lima	lima	0	0	1	0
somrarna	the summers	0	0	1	0
somrarna	summers	0	0	1	0
skivbolag	record label	0	0	1	0
skivbolag	record company	0	0	1	0
framgångsrik	successful	0	0	1	1
kinesisk	chinese	0	0	1	1
skotsk	scottish	0	0	1	1
chi	chi	0	0	1	0
gruppspelet	group stage	0	0	1	0
gruppspelet	groupplay	0	0	1	0
gruppspelet	group play	0	0	1	0
nobel	nobel	0	0	1	0
resten	the rest	0	0	1	0
resten	rest	0	0	1	0
planerade	planeade	0	0	1	0
planerade	planned	0	0	1	0
nytta	useful	0	0	1	0
nytta	good	0	0	1	0
nytta	from	0	0	1	0
geografisk	geographic	0	0	1	1
geografisk	geographical	0	0	1	1
geografisk	spatial	0	0	1	0
titanics	titanic's	0	0	1	0
titanics	titanic	0	0	1	0
konkurrens	competition	0	0	1	1
prinsen	prince	0	0	1	0
prinsen	the prince	0	0	1	0
uppstå	develop	0	0	1	0
uppstå	occur	0	0	1	0
uppstå	arise	0	0	1	1
strider	strides	0	0	1	0
strider	battles	0	0	1	0
strider	conflict	0	0	1	0
öppnat	opened	0	0	1	0
öppnat	opening	0	0	1	0
utropade	exclaimed	0	0	1	0
utropade	cried out	0	0	1	0
bakterier	bacteria	0	0	1	0
avsikten	intention	0	0	1	0
avsikten	purpose	0	0	1	0
iii	iii	0	0	1	0
platsen	the place	0	0	1	0
platsen	place	0	0	1	0
platsen	site	0	0	1	0
ansvaret	responsibility	0	0	1	0
ansvaret	the responsiblity	0	0	1	0
britney	britney	0	0	1	0
f	f	0	0	1	1
tunnel	tunnel	0	0	1	1
gabriel	gabriel	0	0	1	0
baserad	based	0	0	1	1
kedja	chain	0	0	1	1
tillgång	access	0	0	1	0
kategorisvenska	category: swedish	0	0	1	0
direkt	direct	0	0	1	1
direkt	directly	0	0	1	1
baseras	based on	0	0	1	0
baseras	bases	0	0	1	0
baseras	based	0	0	1	0
baserar	base	0	0	1	0
baserar	based	0	0	1	0
bestämde	determined	0	0	1	0
bestämde	chose	0	0	1	0
baserat	based	0	0	1	0
kyrkan	the church	0	0	1	0
kyrkan	church	0	0	1	0
indianerna	the indians	0	0	1	0
indianerna	indians	0	0	1	0
titlar	titles	0	0	1	0
do	do	0	0	1	1
hänvisning	reference	0	0	1	1
allians	alliance	0	0	1	1
konstnärliga	artistic	0	0	1	0
holländska	dutch	0	0	1	1
hållas	be	0	0	1	0
hållas	be held	0	0	1	0
ärkebiskop	archbishop	0	0	1	1
cecilia	cecilia	0	0	1	0
fett	fat	0	0	1	1
democracy	democracy	0	0	1	0
internationellt	international	0	0	1	0
internationellt	internationally	0	0	1	1
tränaren	coach	0	0	1	0
tränaren	the coach	0	0	1	0
tränaren	trans breaker	0	0	1	0
räknade	calculated	0	0	1	0
räknade	counted	0	0	1	0
lanserade	introduced	0	0	1	0
lanserade	launched	0	0	1	0
internationella	international	0	0	1	0
vilhelm	vilhelm	0	0	1	0
fångenskap	captivity	0	0	1	1
revs	described	0	0	1	0
revs	was demolished	0	0	1	0
rousseau	rousseau	0	0	1	0
riktig	real	0	0	1	0
klar	clear	0	0	1	1
klar	done	0	0	1	0
trycktes	was published	0	0	1	0
trycktes	printed	0	0	1	0
fram	until	0	0	1	0
fram	out	0	0	1	1
herrlandskamper	herrlandskamper	0	0	1	0
herrlandskamper	men's international contest	0	0	1	0
herrlandskamper	men's international contests	0	0	1	0
förlaget	publisher	0	0	1	0
förlaget	the publisher	0	0	1	0
förlaget	the publishing company	0	0	1	0
schweiziska	swiss	0	0	1	0
jämnt	even	0	0	1	0
jämnt	evenly	0	0	1	0
gammal	old	0	0	1	1
terrier	terriers	0	0	1	0
terrier	terrier	0	0	1	1
körberg	körberg	0	0	1	0
framträder	stand out	0	0	1	0
framträder	stand	0	0	1	0
framträder	appear	0	0	1	0
dryck	beverage	0	0	1	1
dryck	drink	0	0	1	1
dryck	drinks	0	0	1	0
registrerade	data	0	0	1	0
registrerade	noted	0	0	1	0
överensstämmer	conform	0	0	1	0
överensstämmer	agree	0	0	1	0
överensstämmer	match	0	0	1	0
olyckan	incident	0	0	1	0
olyckan	the accident	0	0	1	0
bilbo	bilbo	0	0	1	0
omslaget	cover	0	0	1	0
omslaget	the cover	0	0	1	0
dy	younger	0	0	1	0
halvklotet	hemisphere	0	0	1	0
strid	conflict	0	0	1	1
strid	fight	0	0	1	1
slöts	concluded	0	0	1	0
slöts	signed	0	0	1	0
industrier	industries	0	0	1	0
le	smile	0	0	1	1
le	le	0	0	1	0
mänskligt	human	0	0	1	0
§	s	0	0	1	0
la	la	0	0	1	1
variationer	variations	0	0	1	0
berget	mount	0	0	1	0
berget	the mountain	0	0	1	0
mänskliga	human	0	0	1	0
lp	lp	0	0	1	0
dess	then	0	0	1	0
dess	its	0	0	1	1
eus	eu	0	0	1	0
träffa	meet	0	0	1	1
träffa	see	0	0	1	1
dag	dag	0	0	1	0
dag	day	0	0	1	1
ägg	agg	0	0	1	0
ägg	eggs	0	0	1	0
ägg	egg	0	0	1	1
spela	play	0	0	1	1
dam	dam	0	0	1	0
dam	lady	0	0	1	1
dan	dan	0	0	1	0
övernaturliga	supernatural	0	0	1	0
övernaturliga	over natural	0	0	1	0
tillkommit	accured	0	0	1	0
tillkommit	been	0	0	1	0
ägs	is owned	0	0	1	0
ägs	(is) owned	0	0	1	0
ägs	owned	0	0	1	0
periodiska	periodic	0	0	1	0
ägt	taken	0	0	1	0
ägt	agt	0	0	1	0
das	das	0	0	1	0
sammanhanget	connection	0	0	1	0
sammanhanget	context	0	0	1	0
guds	god	0	0	1	0
guds	god's	0	0	1	0
day	day	0	0	1	0
kontinuerligt	continuous	0	0	1	0
kontinuerligt	continous	0	0	1	0
utdöda	extinct	0	0	1	0
beslut	decision	0	0	1	1
morris	morris	0	0	1	0
dömdes	sentenced	0	0	1	0
dömdes	was convicted	0	0	1	0
syftade	alluded to	0	0	1	0
syftade	aiming	0	0	1	0
syftade	aimed	0	0	1	0
spridningen	spread	0	0	1	0
spridningen	the spread	0	0	1	0
spridningen	proliferation	0	0	1	0
lysande	brilliant	0	0	1	1
lysande	illuminating	0	0	1	0
förteckning	index	0	0	1	0
förteckning	label	0	0	1	0
förteckning	listing	0	0	1	0
juridisk	legal	0	0	1	1
författarna	the authors	0	0	1	0
författarna	writers	0	0	1	0
emi	emi	0	0	1	0
tillgången	access	0	0	1	0
pitts	pitts	0	0	1	0
kristiansson	kristiansen	0	0	1	0
kristiansson	ristiansson	0	0	1	0
kristiansson	kristiansson	0	0	1	0
företag	company	0	0	1	1
företag	companies	0	0	1	0
företag	business	0	0	1	1
inspirerade	inspired	0	0	1	0
segern	the victory	0	0	1	0
segern	victory	0	0	1	0
marley	marley	0	0	1	0
marley	bob marley = singer	0	0	1	0
arbetskraft	workforce	0	0	1	0
arbetskraft	labor	0	0	1	1
fattigdomen	poverty	0	0	1	0
matt	matt	0	0	1	0
matt	dull	0	0	1	1
jerusalem	jerusalem	0	0	1	1
jamaicanska	jamaican	0	0	1	0
mats	mat's	0	0	1	0
mats	attention	0	0	1	0
intellektuella	intellectuals	0	0	1	0
intellektuella	intellectual	0	0	1	0
ren	deer	0	0	1	0
ren	clean	0	0	1	1
mötley	mötley	0	0	1	0
deras	their	0	0	1	1
red	eds	0	0	1	0
filmatiseringen	film version	0	0	1	0
träning	training	0	0	1	1
träning	practice	0	0	1	1
frank	franks	0	0	1	0
webbplats	website	0	0	1	0
webbplats	site	0	0	1	0
franz	franz	0	0	1	0
odlas	cultured	0	0	1	0
arbetare	workers	0	0	1	0
inleds	starts	0	0	1	0
inleds	start	0	0	1	0
gravid	pregnant	0	0	1	1
referenser	references	0	0	1	0
farbror	uncle	0	0	1	1
inleda	initiate	0	0	1	1
south	south	0	0	1	0
offentlig	public	0	0	1	1
offentlig	published	0	0	1	0
klassisk	classical	0	0	1	1
klassisk	classic	0	0	1	1
färöarna	faroe islands	0	0	1	0
färöarna	the faroe islands	0	0	1	0
pga	because of (short of "på grund av")	0	0	1	0
pga	due	0	0	1	0
uppges	reported	0	0	1	0
uppger	states	0	0	1	0
uppger	state	0	0	1	0
insikt	insight	0	0	1	1
insikt	recognition	0	0	1	0
upphörde	ceased	0	0	1	0
upphörde	expired	0	0	1	0
upphörde	discontinued	0	0	1	0
levnadsstandarden	the standard of living	0	0	1	0
levnadsstandarden	living standard	0	0	1	0
levnadsstandarden	standard of living	0	0	1	0
tillämpa	administer	0	0	1	0
tillämpa	implement	0	0	1	0
tillämpa	applying	0	0	1	0
fruktade	feared	0	0	1	0
veckan	weeks	0	0	1	0
veckan	the week	0	0	1	0
leder	leads	0	0	1	0
leder	leading (to)	0	0	1	0
leder	lead	0	0	1	0
fördrag	agreement	0	0	1	0
fördrag	treaty	0	0	1	1
utlopp	outflow	0	0	1	1
utlopp	outlet	0	0	1	1
kantonerna	the cantons	0	0	1	0
kantonerna	cantons	0	0	1	0
maidens	maidens	0	0	1	0
leden	hinge	0	0	1	0
leden	lines	0	0	1	0
leden	the route	0	0	1	0
palestina	palestine	0	0	1	1
demonstrationer	demonstrations	0	0	1	0
bundna	bonded	0	0	1	0
bundna	tied	0	0	1	0
bundna	bound	0	0	1	0
noterade	note	0	0	1	0
noterade	noted	0	0	1	0
innehade	held	0	0	1	0
innehade	possessed	0	0	1	0
firades	celebrated	0	0	1	0
firades	was	0	0	1	0
firades	was celebrated	0	0	1	0
kvinnlig	females	0	0	1	0
kvinnlig	female	0	0	1	1
bevarats	protected	0	0	1	0
bevarats	preserved	0	0	1	0
läkemedelsverket	food and drug administration	0	0	1	0
läkemedelsverket	medicines work	0	0	1	0
läkemedelsverket	medical products agency	0	0	1	0
domaren	judge	0	0	1	0
domaren	the judge	0	0	1	0
matematisk	mathematical	0	0	1	1
matematisk	mathematic	0	0	1	0
uteslutande	exclusivly	0	0	1	0
uteslutande	only	0	0	1	0
uteslutande	exclusively	0	0	1	1
bröt	brot	0	0	1	0
bröt	broke	0	0	1	0
sweden	sweden	0	0	1	0
kvalificerade	qualifying	0	0	1	0
universum	universe	0	0	1	1
bröd	bread	0	0	1	1
havs	at sea	0	0	1	0
havs	sea	0	0	1	0
aristoteles	aristoteles	0	0	1	0
aristoteles	aristotle	0	0	1	0
tids	time	0	0	1	0
operativsystem	os	0	0	1	0
operativsystem	operative systems	0	0	1	0
operativsystem	operating system	0	0	1	0
basist	bassist	0	0	1	1
have	have	0	0	1	0
idag	today	0	0	1	1
mil	mile	0	0	1	0
mil	swedish miles	0	0	1	0
mil	mil	0	0	1	0
min	my	0	0	1	1
mia	mia	0	0	1	0
erkända	acknowledged	0	0	1	0
erkända	recognized	0	0	1	0
därigenom	by which	0	0	1	0
därigenom	thus	0	0	1	0
därigenom	thereby	0	0	1	1
eget	own	0	0	1	0
kroppar	cells	0	0	1	0
kroppar	bodies	0	0	1	0
tidningar	press	0	0	1	0
tidningar	magazines	0	0	1	0
mig	me	0	0	1	1
mix	mix	0	0	1	1
experter	experts	0	0	1	0
konstverk	work of art	0	0	1	0
konstverk	artworks	0	0	1	0
konstverk	artwork	0	0	1	0
måste	have to	0	0	1	1
måste	must	0	0	1	1
konkurrerande	competing	0	0	1	0
skolgång	school attendance	0	0	1	1
skolgång	schooling	0	0	1	0
resurser	resources	0	0	1	1
resultatet	the result	0	0	1	0
resultatet	result	0	0	1	0
utgörs	consists of	0	0	1	0
utgörs	is	0	0	1	0
utgörs	make up	0	0	1	0
dinosaurier	dinosaurs	0	0	1	0
varandras	each other	0	0	1	0
varandras	each others	0	0	1	0
varandras	each other's	0	0	1	0
befälet	the command	0	0	1	0
befälet	command	0	0	1	0
resultaten	the results	0	0	1	0
resultaten	results	0	0	1	0
epicentrum	epicentre	0	0	1	1
epicentrum	epicenter	0	0	1	1
sist		0	0	1	0
sist	finally	0	0	1	0
sist	last	0	0	1	1
låten	the song	0	0	1	0
låten	song	0	0	1	0
efternamn	last name	0	0	1	1
efternamn	lastname	0	0	1	0
efternamn	surname	0	0	1	1
homogen	homogenous	0	0	1	0
stranden	shore	0	0	1	0
stranden	the beach	0	0	1	0
upprustning	renovation	0	0	1	0
irakkriget	iraq war	0	0	1	0
användare	users	0	0	1	1
republikanska	republican	0	0	1	0
nämns	mentioned	0	0	1	0
upptäckt	discovered	0	0	1	1
upptäckt	found	0	0	1	0
upptäckt	discovery	0	0	1	1
milano	milano	0	0	1	0
upptäcks	discoverd	0	0	1	0
upptäcks	detected	0	0	1	0
upptäcks	is discovered	0	0	1	0
deuterium	deuterium	0	0	1	0
tidskrift	newspaper	0	0	1	0
tidskrift	magazine	0	0	1	1
capita	capita	0	0	1	0
styrke	strength	0	0	1	0
styrke	been	0	0	1	0
upptäcka	detection	0	0	1	0
upptäcka	discover	0	0	1	1
viktigaste	most important	0	0	1	0
styrka	strength	0	0	1	1
styrka	power	0	0	1	1
text	text	0	0	1	1
charles	charles	0	0	1	0
hamlet	hamlet	0	0	1	0
inhemsk	domestic	0	0	1	1
inhemsk	native	0	0	1	1
ugglas	owl	0	0	1	0
ugglas	ugglas	0	0	1	0
igång	start	0	0	1	0
igång	start up	0	0	1	0
fungerade	thought	0	0	1	0
fungerade	working	0	0	1	0
kurfursten	elector	0	0	1	0
sådant	such	0	0	1	0
rytmiska	rhythmic	0	0	1	0
rytmiska	more rhythmic	0	0	1	0
förintelsen	holocaust	0	0	1	0
förintelsen	the genocide	0	0	1	0
sådana	such	0	0	1	0
uganda	uganda	0	0	1	0
temperatur	temperature	0	0	1	1
satan	satan	0	0	1	1
shahen	the shah	0	0	1	0
shahen	shah	0	0	1	0
bryssel	brussels	0	0	1	1
organiska	organic	0	0	1	0
snitt	on average	0	0	1	0
snitt	average	0	0	1	0
arean	the area	0	0	1	0
arean	the space	0	0	1	0
arean	area	0	0	1	0
buddhismen	buddhism	0	0	1	0
buddhismen	buddism	0	0	1	0
buddhismen	buddhismen	0	0	1	0
regimen	regime	0	0	1	0
studenterna	students	0	0	1	0
studenterna	the students	0	0	1	0
richards	richards	0	0	1	0
högskola	college	0	0	1	0
vinsten	the win	0	0	1	0
vinsten	gain	0	0	1	0
organ	body	0	0	1	0
organ	agency	0	0	1	0
organ	organ	0	0	1	1
nazitysklands	nazi germany	0	0	1	0
nazitysklands	nazi germany's	0	0	1	0
angränsande	adjoining	0	0	1	1
angränsande	adjacent	0	0	1	1
vinster	profit	0	0	1	0
vinster	gains	0	0	1	0
majoriteten	the majority	0	0	1	0
lyckade	successful	0	0	1	0
borde	should	0	0	1	1
byggdes	was	0	0	1	0
byggdes	was built	0	0	1	0
möjligheterna	possibilities	0	0	1	0
möjligheterna	the possibilities	0	0	1	0
krävde	demanded	0	0	1	0
ålands	Åland island's	0	0	1	0
ålands	the Åland island's	0	0	1	0
ålands	aland	0	0	1	0
national	national	0	0	1	0
fåglarnas	the birds'	0	0	1	0
fåglarnas	birds	0	0	1	0
svenska	swedish	0	0	1	1
eleonora	eleonora	0	0	1	0
kapitalet	the capital	0	0	1	0
kapitalet	capital	0	0	1	0
svenskt	swedish	0	0	1	0
egentlig	actual; factual; real	0	0	1	0
egentlig	actual	0	0	1	0
bokförlaget	publisher	0	0	1	0
bokförlaget	bokförlaget	0	0	1	0
bokförlaget	publishing house	0	0	1	0
debutalbumet	the debut-album	0	0	1	0
debutalbumet	debut album	0	0	1	0
reform	reform	0	0	1	1
offentligt	public	0	0	1	0
offentligt	publicly	0	0	1	0
konverterade	converted	0	0	1	0
ordnade	arranged	0	0	1	0
ordnade	parent	0	0	1	0
bruno	bruno	0	0	1	0
carlsson	carlsson	0	0	1	0
avslutades	ended; concluded	0	0	1	0
avslutades	closed	0	0	1	0
avslutades	concludes	0	0	1	0
ordentligt	proper	0	0	1	0
ordentligt	properly	0	0	1	1
ordentligt	firmly	0	0	1	0
förekommer	occurs	0	0	1	0
förekommer	preferred is	0	0	1	0
koncept	concept	0	0	1	0
industrialisering	industrialization	0	0	1	1
tobias	tobias	0	0	1	0
uppskattade	estimated	0	0	1	0
uppskattade	appreciated	0	0	1	0
listan	the list	0	0	1	0
viktigare	important	0	0	1	0
viktigare	more important	0	0	1	0
buddhas	buddha's	0	0	1	0
buddhas	buddhas	0	0	1	0
konservativa	conservative	0	0	1	0
övrigt	other	0	0	1	0
miniatyr|karta	thumbnail map	0	0	1	0
miniatyr|karta	miniature|map	0	0	1	0
litteratur	literature	0	0	1	1
litteratur	litterature	0	0	1	0
aktuellt	current	0	0	1	0
aktuellt	relevant	0	0	1	0
kommunicerar	communicates	0	0	1	0
regimer	regimens	0	0	1	0
regimer	regimes	0	0	1	0
aktuella	current	0	0	1	0
sachsen	saxony	0	0	1	1
sachsen	sachsen	0	0	1	0
fester	celebrations	0	0	1	0
fester	parties	0	0	1	0
befolkningstätheten	population density	0	0	1	0
befolkningstätheten	n/a	0	0	1	0
befolkningstätheten	state of the population	0	0	1	0
inneburit	meant	0	0	1	0
inneburit	resulted	0	0	1	0
befogenhet	warrant	0	0	1	0
befogenhet	authority	0	0	1	1
befogenhet	authorization	0	0	1	0
medicinsk	medical	0	0	1	1
elektroner	electron	0	0	1	0
elektroner	electrons	0	0	1	0
news	news	0	0	1	0
kär	carboxyl	0	0	1	0
kär	in love	0	0	1	1
ad	ad	0	0	1	0
tunisien	tunisia	0	0	1	0
grupperingar	grouping	0	0	1	0
grupperingar	groups	0	0	1	0
grupperingar	groupings	0	0	1	0
slippa	avoid	0	0	1	1
gaza	gaza	0	0	1	0
igen	again	0	0	1	1
igen	back	0	0	1	1
igen	recognize	0	0	1	0
döden	death	0	0	1	0
lätta	light	0	0	1	0
lätta	lighten	0	0	1	1
define	define	0	0	1	0
asteroider	astroids	0	0	1	0
asteroider	asteroids	0	0	1	0
samhällen	communities	0	0	1	0
samhällen	societies	0	0	1	0
väljas	elected	0	0	1	0
väljas	be elected	0	0	1	0
väljas	choose	0	0	1	0
stationen	station	0	0	1	0
stationer	stations	0	0	1	0
orange	orange	0	0	1	1
vänsterpartiet	leftist party	0	0	1	0
vänsterpartiet	left-wing party	0	0	1	0
vänsterpartiet	left wing party	0	0	1	0
prestigefyllda	prestigious	0	0	1	0
nederländerna	the netherlands	0	0	1	0
nederländerna	netherlands	0	0	1	1
napoleon	napoleon	0	0	1	1
samhället	the society	0	0	1	0
samhället	society	0	0	1	0
augusti	august	0	0	1	1
bruket	use	0	0	1	0
bruket	the use	0	0	1	0
stalin	stalin	0	0	1	0
ar	is	0	0	1	0
klassificera	classifying	0	0	1	0
klassificera	classify	0	0	1	1
betraktade	considered	0	0	1	0
betraktade	watched	0	0	1	0
när	when	0	0	1	1
externa	external	0	0	1	0
nät	web	0	0	1	1
nät	net(work)	0	0	1	0
palats	palaces	0	0	1	0
palats	palace	0	0	1	1
tagits	taken	0	0	1	0
flyktingar	refugees	0	0	1	0
slöt	joined (in peace)	0	0	1	0
slöt	closed	0	0	1	0
betalade	payed	0	0	1	0
betalade	paid	0	0	1	0
vistelse	visit	0	0	1	1
vistelse	stay	0	0	1	1
nått	reached	0	0	1	0
prosa	prose	0	0	1	1
goebbels	goebbels	0	0	1	0
goebbels	geobbels	0	0	1	0
låg	low	0	0	1	1
administration	administration	0	0	1	1
födda	born	0	0	1	0
fördes	sea were entered	0	0	1	0
fördes	out	0	0	1	0
förhindrar	prevents	0	0	1	0
förhindrar	prevent	0	0	1	0
födde	gave birth too	0	0	1	0
födde	born	0	0	1	0
wolfgang	wolfgang	0	0	1	0
blodtrycket	the blood pressure	0	0	1	0
blodtrycket	blood pressure	0	0	1	0
fler	more	0	0	1	0
hinduismen	hinduism	0	0	1	0
hinduismen	up	0	0	1	0
kallad	known as the	0	0	1	0
kallad	know as	0	0	1	0
kallad	called	0	0	1	1
kontrollera	control	0	0	1	1
kontrollera	controlling	0	0	1	0
torbjörn	torbjörn	0	0	1	0
torbjörn	torbjorn	0	0	1	0
värnpliktiga	conscripted	0	0	1	0
värnpliktiga	inductees	0	0	1	0
kallat	called	0	0	1	0
bönorna	bean	0	0	1	0
bönorna	beans	0	0	1	0
kallas	called	0	0	1	0
vanliga	ordinary	0	0	1	0
vanliga	regular	0	0	1	0
vanliga	usual	0	0	1	1
center	center	0	0	1	1
thailand	thailand	0	0	1	0
seth	seth	0	0	1	0
antonio	antonio	0	0	1	0
sett	seen	0	0	1	1
sett	except	0	0	1	0
hoppas	hope	0	0	1	1
svensk	swedish	0	0	1	1
undvika	prevent	0	0	1	0
undvika	avoid	0	0	1	1
position	position	0	0	1	1
rush	rush	0	0	1	1
isär	ice	0	0	1	0
isär	apart	0	0	1	1
stores	great	0	0	1	0
stores	the great	0	0	1	0
stores	the great's	0	0	1	0
kontaktade	contacted	0	0	1	0
folkrepubliken	people's republic	0	0	1	0
folkrepubliken	people"s republic	0	0	1	0
mystiska	mysterious	0	0	1	0
mystiska	mystical	0	0	1	0
mystiska	mysiska	0	0	1	0
wagner	wagner	0	0	1	0
grekiskans	the greek's	0	0	1	0
grekiskans	greek	0	0	1	0
flertal	several	0	0	1	0
flertal	majority group	0	0	1	0
vanligt	normal	0	0	1	0
vanligt	usual	0	0	1	0
kampf	on	0	0	1	0
kampf	kampf	0	0	1	0
liverpools	liverpool's	0	0	1	0
liverpools	liverpools	0	0	1	0
reformer	reformers	0	0	1	0
reformer	reforms	0	0	1	0
lake	lake	0	0	1	0
mentala	mental	0	0	1	0
mentala	mentala	0	0	1	0
underhållning	entertainment	0	0	1	1
huvudstäder	capital cities	0	0	1	0
huvudstäder	capitals	0	0	1	0
streck	bar	0	0	1	0
belgrad	belgrade	0	0	1	1
läsare	reader	0	0	1	1
läsare	readers	0	0	1	0
lika	similar	0	0	1	1
lika	alike	0	0	1	1
lika	equal	0	0	1	1
dubai	dubai	0	0	1	0
jämför	compare	0	0	1	0
koden	the code	0	0	1	0
koden	code	0	0	1	0
användningen	use	0	0	1	0
användningen	the use	0	0	1	0
chrusjtjov	khrushchev	0	0	1	0
chrusjtjov	chrusjtjov	0	0	1	0
höger	right	0	0	1	1
höger	hoger	0	0	1	0
likt	like	0	0	1	1
kejsarens	emperor	0	0	1	0
kejsarens	the emperor's	0	0	1	0
kejsarens	emperors	0	0	1	0
works	works	0	0	1	0
släpper	release	0	0	1	0
släpper	releases	0	0	1	0
albumets	album	0	0	1	0
albumets	album's	0	0	1	0
albumets	albuments	0	0	1	0
starkaste	strongest	0	0	1	0
starkaste	the strongest	0	0	1	0
dvärgar	dwarves	0	0	1	0
dvärgar	dwarfs	0	0	1	0
känsla	feeling	0	0	1	1
känsla	sense	0	0	1	1
insats	contribution	0	0	1	1
insats	intermediate	0	0	1	0
insats	stake	0	0	1	1
etablerades	established	0	0	1	0
etablerades	was established	0	0	1	0
minsta	minimum	0	0	1	0
dött	died	0	0	1	0
dött	dead	0	0	1	0
dött	dott	0	0	1	0
ungarna	the kids	0	0	1	0
ungarna	kids	0	0	1	0
ungarna	the young	0	0	1	0
est	est	0	0	1	0
gänget	the group	0	0	1	0
gänget	the gang	0	0	1	0
gänget	gang	0	0	1	0
joachim	joachim	0	0	1	0
påminde	reminded	0	0	1	0
skildrar	describes	0	0	1	0
skildrar	depicts	0	0	1	0
skildrar	portrays	0	0	1	0
kategorifiktiva	category fictitious	0	0	1	0
gisslan	hostage	0	0	1	1
gisslan	hostages	0	0	1	0
hjärnan	brain	0	0	1	0
hjärnan	the brain	0	0	1	0
internationalen	international	0	0	1	0
definitionen	definition	0	0	1	0
definitionen	the definition	0	0	1	0
nattetid	overnight	0	0	1	0
definitioner	definitions	0	0	1	0
mjölk	milk	0	0	1	1
säkerhetsrådet	security	0	0	1	0
starkare	strong	0	0	1	0
starkare	stronger	0	0	1	0
leopold	leopold	0	0	1	0
förklaring	explaination	0	0	1	0
förklaring	explanation	0	0	1	1
förklaring	statement	0	0	1	0
nordkorea	north korea	0	0	1	0
nordkorea	north koreans	0	0	1	0
socker	sugar	0	0	1	1
glada	happy	0	0	1	0
tomt	empty	0	0	1	0
tomt	blank	0	0	1	0
andel	percentage	0	0	1	0
andel	share	0	0	1	1
anden	the holy spirit	0	0	1	0
anden	spirit	0	0	1	0
alexanders	alexanders	0	0	1	0
alexanders	alexander's	0	0	1	0
kapital	capital	0	0	1	1
omgiven	surrounded	0	0	1	1
potatis	potato	0	0	1	1
växter	plants	0	0	1	0
mått	measurements	0	0	1	0
mått	measure	0	0	1	1
mått	measurement	0	0	1	1
monarken	the monarch	0	0	1	0
monarken	monarch	0	0	1	0
chris	chris	0	0	1	0
rösta	vote	0	0	1	1
nordsjön	north sea	0	0	1	1
ljusare	brighter	0	0	1	0
ljusare	lighter	0	0	1	0
vimmerby	vimmerby	0	0	1	0
hatar	hate	0	0	1	0
hatar	hates	0	0	1	0
ridge	ridge	0	0	1	0
densamma	the same	0	0	1	0
densamma	same	0	0	1	0
försvara	research be	0	0	1	0
försvara	defend	0	0	1	1
försvara	defending	0	0	1	0
avrättades	was executed	0	0	1	0
avrättades	executed	0	0	1	0
illuminati	illuminati	0	0	1	0
västerut	west	0	0	1	1
västerut	westward; west	0	0	1	0
västerut	westwards	0	0	1	0
kuben	cube	0	0	1	0
kuben	the cube	0	0	1	0
tronföljare	heir	0	0	1	0
tronföljare	heir apparent	0	0	1	0
tronföljare	successor	0	0	1	0
flyg	flight	0	0	1	0
flyg	airforce	0	0	1	0
flyg	air	0	0	1	0
klockan	o'clock	0	0	1	1
klockan	clock	0	0	1	0
civilbefolkningen	civilian population	0	0	1	0
civilbefolkningen	the civilian population	0	0	1	0
civilbefolkningen	civilians	0	0	1	0
ryssarna	the russians	0	0	1	0
ryssarna	russians	0	0	1	0
brand	fire	0	0	1	1
ättlingar	descendants	0	0	1	0
flygvapnet	air force	0	0	1	0
flygvapnet	the airforce	0	0	1	0
kraft	force	0	0	1	1
kraft	power	0	0	1	1
bud	bid	0	0	1	1
bud	bids	0	0	1	0
bud	message	0	0	1	1
årtionden	decades	0	0	1	0
utsåg	declared	0	0	1	0
utsåg	appointed	0	0	1	0
vetenskap	science	0	0	1	1
utrymme	space	0	0	1	1
västra	west	0	0	1	1
västra	vastra	0	0	1	0
västra	western	0	0	1	1
lissabon	lissabon	0	0	1	0
lissabon	lisbon	0	0	1	1
australiens	australia	0	0	1	0
australiens	australia's	0	0	1	0
kuiperbältet	the cuyper belt	0	0	1	0
kuiperbältet	kuiperbaltet	0	0	1	0
kuiperbältet	the kuiper belt	0	0	1	0
nedre	lower	0	0	1	1
nedre	bottom	0	0	1	0
kaffe	coffee	0	0	1	1
minuter	minutes	0	0	1	1
täcker	attacks	0	0	1	0
täcker	covers	0	0	1	0
circus	circus	0	0	1	0
paraguay	paraguay	0	0	1	1
tolkningen	interpretetation	0	0	1	0
tolkningen	interpretation	0	0	1	0
omloppsbanor	orbits	0	0	1	0
omloppsbanor	orbit	0	0	1	0
anhöriga	relatives	0	0	1	0
anhöriga	kin	0	0	1	0
autism	autism	0	0	1	1
skador	damage	0	0	1	0
manlig	male	0	0	1	1
manlig	manly	0	0	1	1
identitet	identity	0	0	1	1
besläktade	related	0	0	1	0
proteiner	proteins	0	0	1	0
einsteins	einstein	0	0	1	0
einsteins	once a	0	0	1	0
einsteins	einsteins	0	0	1	0
sandy	sandy	0	0	1	0
gränserna	borders	0	0	1	0
gränserna	the borders	0	0	1	0
gränserna	limits	0	0	1	0
picchu	picchu	0	0	1	0
stimulans	stimulation	0	0	1	1
stimulans	stimulating	0	0	1	0
betonade	emphasized	0	0	1	0
endast	only	0	0	1	1
endast	merely	0	0	1	1
uppfatta	apprehend	0	0	1	1
uppfatta	perceived	0	0	1	0
uppfatta	perceive	0	0	1	1
astronomi	astronomy	0	0	1	1
variation	diversity	0	0	1	0
variation	variety	0	0	1	1
akademisk	academical	0	0	1	1
akademisk	academic	0	0	1	1
cirkel	circular	0	0	1	0
föräldrarna	the parents	0	0	1	0
föräldrarna	parents	0	0	1	0
föräldrarna	foraldrama	0	0	1	0
philips	philips	0	0	1	0
fakta	facts	0	0	1	0
fakta	fact	0	0	1	0
inträde	entry	0	0	1	1
attacker	attacks	0	0	1	0
attacker	assaults	0	0	1	0
baker	baker	0	0	1	0
baker	panadero	0	0	1	0
svag	weak	0	0	1	1
uppfattningen	comprehension	0	0	1	0
uppfattningen	view	0	0	1	0
fönster	windows	0	0	1	0
fönster	window	0	0	1	1
återställa	reset	0	0	1	1
återställa	restore	0	0	1	1
återställa	resett	0	0	1	0
stämma	stutter	0	0	1	0
stämma	sue	0	0	1	1
stämma	meeting	0	0	1	1
ögon	eye (-s)	0	0	1	0
ögon	eyes	0	0	1	0
nelson	nelson	0	0	1	1
brottslingar	criminals	0	0	1	0
förespråkare	spokesman	0	0	1	0
förespråkare	proponent	0	0	1	0
slogs	fought	0	0	1	0
slogs	was	0	0	1	0
kännetecknas	characterized (by)	0	0	1	0
kännetecknas	is characterized	0	0	1	0
kännetecknas	characterized	0	0	1	0
arkitekt	architect	0	0	1	1
antisemitiska	antisemetic	0	0	1	0
antisemitiska	anti-semitic	0	0	1	0
antisemitiska	antisemitic	0	0	1	0
ozzy	ozzy	0	0	1	0
granskning	review	0	0	1	0
anfallet	the attack	0	0	1	0
anfallet	attack	0	0	1	0
islamisk	islamic	0	0	1	1
paris	paris	0	0	1	1
deltagit	part	0	0	1	0
deltagit	participated	0	0	1	0
tillräckligt	sufficient	0	0	1	0
linköping	linköping	0	0	1	0
kapacitet	the capacity	0	0	1	0
kapacitet	capacity	0	0	1	1
under	during	0	0	1	1
under	for	0	0	1	1
under	under	0	0	1	1
nordost	north east	0	0	1	0
nordost	northeast	0	0	1	0
nordost	the northeast	0	0	1	0
pommern	pommern	0	0	1	0
pommern	pomerania	0	0	1	0
tillåtna	allowed	0	0	1	0
tjänar	earns	0	0	1	0
tjänar	serves	0	0	1	0
förstås	course	0	0	1	0
förstås	mean:	0	0	1	0
förstår	understand	0	0	1	0
förstår	forstar	0	0	1	0
jack	jack	0	0	1	1
evert	everted	0	0	1	0
evert	evert	0	0	1	0
myntade	coined	0	0	1	0
längre	longer	0	0	1	0
tagit	taken	0	0	1	0
tagit	received	0	0	1	0
school	school	0	0	1	0
plural	plural	0	0	1	0
trettioåriga	13 year olds	0	0	1	0
trettioåriga	thirty year's (war)	0	0	1	0
trettioåriga	thirty years	0	0	1	0
venus	venus	0	0	1	1
petersburg	petersburg	0	0	1	0
matematik	mathematic	0	0	1	0
matematik	mathematics	0	0	1	1
verklig	real	0	0	1	1
reklam	advertising	0	0	1	1
reklam	advertisement	0	0	1	1
parten	party	0	0	1	0
ingripande	negative	0	0	1	0
ingripande	intervention	0	0	1	1
rätta	correct	0	0	1	1
rätta	come to grips; court; correct	0	0	1	0
street	street	0	0	1	0
parter	party	0	0	1	0
parter	sides	0	0	1	0
manus	script	0	0	1	1
indierna	the indians	0	0	1	0
indierna	indians	0	0	1	0
stridigheter	oppositions	0	0	1	0
stridigheter	strife	0	0	1	0
aktivt	active	0	0	1	0
aktivt	actively	0	0	1	0
drivande	drive	0	0	1	0
drivande	driving	0	0	1	1
ebba	die	0	0	1	0
ebba	ebba	0	0	1	0
notera	note	0	0	1	1
liberty	liberty	0	0	1	0
journalist	journalist	0	0	1	1
aktiva	active	0	0	1	0
zink	zinc	0	0	1	1
följande	following	0	0	1	1
följande	the following	0	0	1	0
genomföras	carried out	0	0	1	0
genomföras	be performed	0	0	1	0
genomföras	carry out	0	0	1	0
kub	cube	0	0	1	1
disney	disney	0	0	1	0
egyptens	egypt	0	0	1	0
egyptens	egypts	0	0	1	0
egyptens	egypt's	0	0	1	0
zach	zach	0	0	1	0
prata	talk	0	0	1	1
hjälpte	helped	0	0	1	0
flera	many	0	0	1	1
flera	multiple	0	0	1	0
medelhavsklimat	mediterranean climate	0	0	1	0
utredning	study	0	0	1	0
utredning	investigation	0	0	1	1
beck	beck	0	0	1	0
beck	pitch	0	0	1	1
parlamentariska	parliamentary	0	0	1	0
parlamentariska	the parliamentary	0	0	1	0
preparat	substance	0	0	1	0
preparat	preparations	0	0	1	0
preparat	compound	0	0	1	0
studio	studio	0	0	1	1
rysk	russian	0	0	1	1
församling	congregation	0	0	1	1
församling	assembly	0	0	1	1
fördelade	divided	0	0	1	0
fördelade	distributed	0	0	1	0
komplex	complex	0	0	1	1
komplex	komplex	0	0	1	0
studie	study	0	0	1	1
övervägande	the predominant	0	0	1	0
övervägande	predominant	0	0	1	1
övervägande	predominantly	0	0	1	0
forum	forum	0	0	1	1
lagras	stored	0	0	1	0
ty	for	0	0	1	1
giftsnokar	elapidaes	1	0	1	0
giftsnokar	venomous conks	1	0	1	0
giftsnokar	venomous grass snake	1	0	1	0
giftsnokar	passed	1	0	1	0
giftsnokar	venomous snakes	1	0	1	0
giftsnokar	elapidae	1	1	0	0
giftsnokar	elipidae	1	0	1	0
giftsnokar	poisonous snakes	1	1	0	0
giftsnokar	giftsnoakar	1	0	1	0
giftsnokar	venomous snake	1	0	1	0
giftsnokar	elapids	1	1	0	0
giftsnokar	venom	1	0	1	0
giftsnokar	located	1	0	1	0
giftsnokar	poison snakes	1	0	1	0
giftsnokar	toxic snooping	1	0	1	0
giftsnokar	venom snooping	1	0	1	0
precis	precisely	0	0	1	1
precis	just	0	0	1	1
precis	exactly; precisely	0	0	1	0
proportioner	proportions	0	0	1	0
svante	svante	0	0	1	0
isen	the ice	0	0	1	0
kväve	kave	0	0	1	0
kväve	nitrogen	0	0	1	1
strax	soon	0	0	1	0
strax	just	0	0	1	1
julie	julie	0	0	1	0
erektion	erection	0	0	1	1
julia	julia	0	0	1	0
nazistiska	nazi	0	0	1	0
hittades	was found	0	0	1	0
misslyckats	failed	0	0	1	0
volym	volume	0	0	1	1
mattias	mattias	0	0	1	0
klassas	classified	0	0	1	0
vinst	profit	0	0	1	1
vinst	win	0	0	1	1
miniatyr|px|en	miniature	0	0	1	0
konserterna	the concerts	0	0	1	0
konserterna	concerts	0	0	1	0
skicka	send	0	0	1	1
väckte	awakened	0	0	1	0
väckte	aroused	0	0	1	0
behandlingar	treatments	0	0	1	0
samhälle	society	0	0	1	1
södra	southern	0	0	1	0
södra	south	0	0	1	0
inför	before	0	0	1	1
förändringar	changes	0	0	1	0
erhöll	obtained	0	0	1	0
erhöll	recieved	0	0	1	0
erhöll	acquire	0	0	1	0
muse	muse	0	0	1	0
ludvig	louis	0	0	1	0
ludvig	ludvig	0	0	1	0
råkar	happens	0	0	1	0
råkar	happens to	0	0	1	0
vagnar	carts	0	0	1	0
vagnar	wagons	0	0	1	0
vagnar	carriges	0	0	1	0
fermentering	fermentation	0	0	1	0
avsätta	unseat	0	0	1	1
avsätta	depositing	0	0	1	0
belgiens	belgium	0	0	1	0
belgiens	belgium's	0	0	1	0
igelkottens	the hedgehog's	0	0	1	0
igelkottens	hedgehog	0	0	1	0
ämne	substance	0	0	1	1
ämne	subject	0	0	1	1
henri	henri - it's a name	0	0	1	0
henri	henri	0	0	1	0
mm	millimeter	0	0	1	0
mm	etc.	0	0	1	0
lukas	luke	0	0	1	1
lukas	lukas	0	0	1	0
antiken	the ancient world	0	0	1	0
antiken	antiquity	0	0	1	0
ms	motor ship	0	0	1	0
henry	henry	0	0	1	1
johanssons	johanssons	0	0	1	0
johanssons	johansson	0	0	1	0
ernest	ernest	0	0	1	0
utgick	started	0	0	1	0
utgick	was deleted	0	0	1	0
partiets	the party's	0	0	1	0
partiets	parties	0	0	1	0
hämtar	download	0	0	1	0
hämtar	is	0	0	1	0
hämtar	gets	0	0	1	0
västerås	västerås	0	0	1	0
västerås	vasteras	0	0	1	0
värvade	recruited	0	0	1	0
värvade	referred	0	0	1	0
persien	persia	0	0	1	0
florida	florida	0	0	1	1
belägna	located	0	0	1	0
belägna	disposed	0	0	1	0
ätten	the dynasty	0	0	1	0
ätten	ater	0	0	1	0
ätten	dynasty	0	0	1	0
ena	one	0	0	1	1
end	end	0	0	1	0
eng	eng.	0	0	1	0
eng	eng	0	0	1	0
iiis	iii's	0	0	1	0
iiis	3's	0	0	1	0
ens	even	0	0	1	0
ens	one's	0	0	1	0
gata	street	0	0	1	1
rörlighet	movement	0	0	1	0
rörlighet	mobility	0	0	1	1
elektriskt	electric	0	0	1	0
elizabeth	elizabeth	0	0	1	0
beskrev	depicted	0	0	1	0
beskrev	described	0	0	1	0
mest	most	0	0	1	1
mest	mostly	0	0	1	1
miniatyr|px|ett	miniature	0	0	1	0
väster	west	0	0	1	1
elektriska	electrical	0	0	1	0
omgångar	in turns; periods; mandates	0	0	1	0
omgångar	cycles	0	0	1	0
åsikt	opinion	0	0	1	1
må	feel	0	0	1	1
må	may	0	0	1	1
må	mon	0	0	1	0
nagasaki	nagasaki	0	0	1	0
kategorier	categories	0	0	1	0
kubanska	cuban	0	0	1	0
tsar	tsar	0	0	1	1
tsar	czar	0	0	1	1
galilei	galilei	0	0	1	0
beteenden	behavior	0	0	1	0
kontrollen	control	0	0	1	0
kontrollen	the control	0	0	1	0
existera	exist	0	0	1	1
beskrivit	described	0	0	1	0
partierna	political parties	0	0	1	0
partierna	portions	0	0	1	0
arbetar	work	0	0	1	0
arbetar	works	0	0	1	0
kejsare	emperor	0	0	1	1
ledamöterna	the commissioners	0	0	1	0
ledamöterna	commisioners	0	0	1	0
ledamöterna	the members	0	0	1	0
kampen	the fight	0	0	1	0
kampen	the struggle	0	0	1	0
kampen	fight	0	0	1	0
over	over	0	0	1	1
fall	where	0	0	1	0
arresterades	was arrested	0	0	1	0
vitt	white	0	0	1	1
vitt	widely	0	0	1	1
london	london	0	0	1	1
synonymt	synonymous	0	0	1	0
synonymt	synonymously	0	0	1	0
frivillig	optional	0	0	1	1
vita	white	0	0	1	1
expansion	expansion	0	0	1	1
bibelns	the bibel's	0	0	1	0
bibelns	the bible's	0	0	1	0
bibelns	bible	0	0	1	0
brinner	on fire	0	0	1	0
brinner	burns	0	0	1	0
brinner	burn	0	0	1	0
ursprungsbefolkningen	the native population	0	0	1	0
ursprungsbefolkningen	indigenous people	0	0	1	0
ursprungsbefolkningen	indigenous population	0	0	1	0
imf	imf	0	0	1	0
edith	edith	0	0	1	0
träd	into	0	0	1	0
träd	tree	0	0	1	1
nytt	new	0	0	1	0
statschef	head of state	0	0	1	0
först	first	0	0	1	1
blott	merely	0	0	1	1
blott	only	0	0	1	1
blott	mere	0	0	1	1
historiens	historys	0	0	1	0
historiens	history's	0	0	1	0
dem	those	0	0	1	1
senast	last (time)	0	0	1	0
senast	last	0	0	1	1
mål	case	0	0	1	1
mål	goal	0	0	1	1
mål	mal	0	0	1	0
produktion	production	0	0	1	1
upptagen	included	0	0	1	0
upptagen	busy	0	0	1	1
upptagen	occupied	0	0	1	1
lämplig	suitable	0	0	1	1
avskaffandet	elimination	0	0	1	0
avskaffandet	abolition	0	0	1	0
avskaffandet	abolishment	0	0	1	0
ansvarar	charge	0	0	1	0
ansvarar	responsible	0	0	1	0
alex	alex	0	0	1	0
miljoner	milions	0	0	1	0
miljoner	millon	0	0	1	0
miljoner	one million	0	0	1	0
miljoner	millions	0	0	1	0
detroit	detroit	0	0	1	0
bunny	bunny	0	0	1	0
sauron	sauron	0	0	1	0
newport	newport	0	0	1	0
storlek	size	0	0	1	1
ursprungligen	initially	0	0	1	0
ursprungligen	originally	0	0	1	1
gälla	valid	0	0	1	0
gälla	be valid	0	0	1	1
äventyr	adventure	0	0	1	1
äventyr	adventures	0	0	1	0
gymnasium	high school	0	0	1	0
bra	good	0	0	1	1
sångaren	singer	0	0	1	0
sångaren	the singer	0	0	1	0
raid	raid	0	0	1	0
förebild	model	0	0	1	1
förebild	role model	0	0	1	0
påtagligt	substantially	0	0	1	0
påtagligt	considerably	0	0	1	0
påtagligt	markedly	0	0	1	0
nio	nine	0	0	1	1
gom	palate	1	1	0	1
gom	corresponding	1	0	1	0
gom	gum	1	0	1	0
gom	mouth	1	1	0	0
gom	related	1	0	1	0
gom	roof of mouth	1	1	0	0
gom	market organization	1	0	1	0
god	good	0	0	1	1
receptorer	receptors	0	0	1	0
ammoniak	ammonia	0	0	1	1
hemland	homeland	0	0	1	1
riktning	direction	0	0	1	1
danmarks	denmarks	0	0	1	0
danmarks	denmark's	0	0	1	0
paulus	paulus	0	0	1	0
paulus	paul	0	0	1	0
got	got	0	0	1	0
independence	independence	0	0	1	0
sätts	is	0	0	1	0
sätts	turned (on)	0	0	1	0
sätts	is placed	0	0	1	0
icke	non	0	0	1	0
icke	none	0	0	1	1
benämnas	named	0	0	1	0
benämnas	entitle	0	0	1	0
benämnas	entitled	0	0	1	0
herman	herman	0	0	1	0
free	free	0	0	1	0
fred	peace	0	0	1	1
prägel	character	0	0	1	0
prägel	mark	0	0	1	0
sätta	insert	0	0	1	0
sätta	set	0	0	1	1
samlade	collected	0	0	1	0
inom	within	0	0	1	1
inom	in	0	0	1	1
drygt	slightly more than	0	0	1	0
drygt	good	0	0	1	0
drygt	approximately	0	0	1	0
växterna	plants	0	0	1	0
statsministern	the prime minister	0	0	1	0
statsministern	prime minister	0	0	1	0
statsministern	head of state	0	0	1	0
räddade	saved	0	0	1	0
studera	study	0	0	1	1
tolerans	tolerance	0	0	1	1
bredvid	beside	0	0	1	1
bredvid	next to	0	0	1	1
vetenskapliga	scientific	0	0	1	0
godkändes	was approved	0	0	1	0
godkändes	approved	0	0	1	0
befolkade	inhabitated	0	0	1	0
befolkade	populated	0	0	1	0
berättelser	tales	0	0	1	0
berättelser	stories	0	0	1	0
vetenskapligt	scientifically	0	0	1	1
vetenskapligt	scientific	0	0	1	0
transporterar	carrying	0	0	1	0
transporterar	transports	0	0	1	0
transporteras	is transported	0	0	1	0
transporteras	transported	0	0	1	0
nyheter	news	0	0	1	0
atmosfär	atmosphere	0	0	1	1
atmosfär	atmospheric	0	0	1	0
museet	the museum	0	0	1	0
museet	museum	0	0	1	0
museer	museums	0	0	1	0
museer	musser	0	0	1	0
tidigt	early	0	0	1	1
tidigt	at an early stage	0	0	1	0
nhl	nhl	0	0	1	0
institutioner	institutions	0	0	1	0
rikaste	the richest	0	0	1	0
rikaste	richest	0	0	1	0
sexuellt	sexual	0	0	1	0
besökare	visitors	0	0	1	0
militär	military	0	0	1	1
sexuella	sexual	0	0	1	0
nyheten	news	0	0	1	0
mercury	mercury	0	0	1	0
uppgörelse	settlement	0	0	1	1
uppgörelse	agreement	0	0	1	1
uppgörelse	deal	0	0	1	0
utsågs	was	0	0	1	0
utsågs	appointed	0	0	1	0
utsågs	was appointed	0	0	1	0
toy	toy	0	0	1	0
tor	thu	0	0	1	0
tor	thor	0	0	1	1
punkten	the point	0	0	1	0
punkten	point	0	0	1	0
dalar	valleys	0	0	1	0
konventionen	the convention	0	0	1	0
konventionen	convention	0	0	1	0
merkurius	mercury	0	0	1	0
konventioner	conventions	0	0	1	0
ton	tonne	0	0	1	0
ton	tone	0	0	1	1
punkter	points	0	0	1	0
punkter	seq	0	0	1	0
tom	tom	0	0	1	0
uppkommit	generated	0	0	1	0
uppkommit	arisen	0	0	1	0
tog	was	0	0	1	0
tog	took	0	0	1	0
adjektiv	adjective	0	0	1	1
adjektiv	adjectives	0	0	1	0
likaså	also	0	0	1	1
likaså	as well	0	0	1	1
födseln	birth	0	0	1	0
födseln	the birth	0	0	1	0
århundradena	ahundradena	0	0	1	0
århundradena	centuries	0	0	1	0
förfäder	ancestors	0	0	1	0
livealbum	live album	0	0	1	0
skildes	separated	0	0	1	0
skildes	was seperated	0	0	1	0
meddelande	message	0	0	1	1
västkusten	the west coast	0	0	1	0
västkusten	west coast	0	0	1	0
åring	year old	0	0	1	0
åring	years	0	0	1	0
båda	both	0	0	1	1
båda	bath	0	0	1	0
kulturarv	culture heritage	0	0	1	0
kulturarv	cultureheritage	0	0	1	0
kulturarv	cultural heritage	0	0	1	0
territoriella	territorial	0	0	1	0
både	both	0	0	1	1
dramer	dramas	0	0	1	0
dramer	plays	0	0	1	0
slutsats	conclusion	0	0	1	1
uppmuntrade	encouragement	0	0	1	0
uppmuntrade	encouraged	0	0	1	0
nödvändigtvis	by necessity	0	0	1	0
nödvändigtvis	necessarily	0	0	1	1
framförallt	above all	0	0	1	0
framförallt	in particular; above all	0	0	1	0
begär	requests	0	0	1	0
begär	request	0	0	1	0
mördad	murdered	0	0	1	0
mördad	murderd	0	0	1	0
religiöst	religious	0	0	1	0
bridge	bridge	0	0	1	1
rad	range	0	0	1	1
rad	line	0	0	1	1
valde	crowned	0	0	1	0
valde	selected	0	0	1	0
valde	chose	0	0	1	0
flyttades	moved	0	0	1	0
pass	an	0	0	1	0
rak	straight	0	0	1	1
rak	linear	0	0	1	0
sköt	forwarder	0	0	1	0
sköt	shot	0	0	1	0
ras	race	0	0	1	1
ras	ras	0	0	1	0
adhd	adhd	0	0	1	0
åstadkomma	provide	0	0	1	0
åstadkomma	create	0	0	1	1
åstadkomma	achieve	0	0	1	1
tycks	appears	0	0	1	0
ray	ray	0	0	1	0
industriellt	industrially	0	0	1	0
industriellt	industrial	0	0	1	0
hittats	found	0	0	1	0
befruktning	judaism	1	0	1	0
befruktning	fertilization	1	1	0	1
befruktning	conception	1	0	1	1
befruktning	fertilizing	1	0	1	0
befruktning	stimulation	1	0	1	1
befruktning	conceptions	1	0	1	0
befruktning	befrukning	1	0	1	0
befruktning	fertilisation	1	1	0	0
befruktning	insemination	1	1	0	0
befruktning	impregnation	1	1	0	1
befruktning	monograph	1	0	1	0
situationer	situations	0	0	1	0
jorden	the earth	0	0	1	0
jorden	earth	0	0	1	0
jorden	earth; earth; underground	0	0	1	0
lanseringen	the release	0	0	1	0
lanseringen	launch	0	0	1	0
nilsson	nilsson	0	0	1	0
fartyg	vessel	0	0	1	1
fartyg	ship; vessel	0	0	1	0
fartyg	ship	0	0	1	1
industriella	industrial	0	0	1	0
academy	academy	0	0	1	0
situationen	situation	0	0	1	0
situationen	the situation	0	0	1	0
mekaniska	mechanical	0	0	1	0
grundskolan	elementary school	0	0	1	0
tvingas	forced	0	0	1	0
tvingas	system	0	0	1	0
skepp	vessel	0	0	1	1
skepp	ship	0	0	1	1
kärna	core	0	0	1	1
kärna	quarks	0	0	1	0
elektricitet	electricity	0	0	1	1
fralagen	fra law	0	0	1	0
fralagen	fralegen	0	0	1	0
fralagen	the fra law	0	0	1	0
spelat	played	0	0	1	0
spelas	played	0	0	1	0
tanzania	tanzania	0	0	1	0
språken	languages	0	0	1	0
språken	park	0	0	1	0
metal	metal	0	0	1	0
sekt	sect	0	0	1	1
metan	methane	0	0	1	1
språket	language	0	0	1	0
inflytande	influence	0	0	1	1
inflytande	power	0	0	1	0
agnes	agnes	0	0	1	0
utkanten	the outskirts	0	0	1	0
utkanten	outskirts	0	0	1	0
delen	part	0	0	1	0
idrott	sport	0	0	1	1
idrott	sports	0	0	1	1
saga	saga	0	0	1	1
saga	story	0	0	1	0
queen	drottning	0	0	1	0
radio	radio	0	0	1	1
användande	use	0	0	1	0
användande	use; usage	0	0	1	0
förklarade	explained	0	0	1	0
förklarade	said	0	0	1	0
earth	earth	0	0	1	0
sagt	said	0	0	1	0
sagt	i have said	0	0	1	0
radie	radius	0	0	1	1
absolut	absolute; total	0	0	1	0
absolut	absolute	0	0	1	1
skada	damage	0	0	1	1
claude	claude	0	0	1	0
florens	florens	0	0	1	0
florens	florence	0	0	1	1
vinna	win	0	0	1	1
institution	institution	0	0	1	1
gods	domain	0	0	1	0
gods	goods	0	0	1	1
abu	abu	0	0	1	0
andras	others	0	0	1	0
definierat	defined	0	0	1	0
bostadsområden	residential	0	0	1	0
bostadsområden	housing	0	0	1	0
bostadsområden	residential areas	0	0	1	0
nära	close	0	0	1	1
nära	near	0	0	1	1
kommunisterna	communists	0	0	1	0
kommunisterna	communist	0	0	1	0
kommunisterna	the communists	0	0	1	0
guatemala	guatemala	0	0	1	1
präglades	was marked	0	0	1	0
präglades	imprinted	0	0	1	0
präglades	marked	0	0	1	0
gogh	gogh	0	0	1	0
tillhörande	associated	0	0	1	0
tillhörande	belonging to	0	0	1	0
tillhörande	belonging (to)	0	0	1	0
haiti	haiti	0	0	1	1
läsaren	the reader	0	0	1	0
läsaren	reader	0	0	1	0
slags	kind	0	0	1	0
slags	type	0	0	1	0
bläckpenna	statistics	1	0	1	0
bläckpenna	ink pen	1	0	1	0
bläckpenna	ball point pen	1	0	1	0
bläckpenna	pen	1	1	0	0
bläckpenna	ink	1	0	1	0
bläckpenna	ball point pen; pen	1	0	1	0
bläckpenna	balck pen	1	0	1	0
bläckpenna	black pen	1	0	1	0
bläckpenna	quill	1	1	0	0
dödligheten	mortality	0	0	1	0
taubes	taubes	0	0	1	0
kraftiga	strong	0	0	1	0
kraftiga	powerful	0	0	1	0
lovat	promised	0	0	1	0
publicerades	published	0	0	1	0
uppvärmningen	the warmup	0	0	1	0
uppvärmningen	heating	0	0	1	0
uppvärmningen	the warm-up	0	0	1	0
tidningen	the newspaper	0	0	1	0
tidningen	journal	0	0	1	0
tidningen	paper	0	0	1	0
uppsättning	equipment	0	0	1	1
uppsättning	set	0	0	1	1
uppsättning	set of	0	0	1	0
kroppen	body	0	0	1	0
kroppen	the body	0	0	1	0
hämtade	taken	0	0	1	0
hämtade	brought	0	0	1	0
sakta	slowly	0	0	1	1
erkände	confession	0	0	1	0
erkände	acknowledged	0	0	1	0
förts	brought	0	0	1	0
förts	cont	0	0	1	0
ockuperat	occupied	0	0	1	0
kristendomen	chritianity	0	0	1	0
kristendomen	christianity	0	0	1	0
utformade	formed	0	0	1	0
utformade	designed	0	0	1	0
används	use	0	0	1	0
används	used	0	0	1	0
långa	langa	0	0	1	0
långa	long	0	0	1	0
mur	wall	0	0	1	1
indoeuropeiska	indo-european	0	0	1	0
indoeuropeiska	european	0	0	1	0
brinnande	burning	0	0	1	1
antikens	the ancient's	0	0	1	0
antikens	ancient	0	0	1	0
långt	far	0	0	1	1
långt	long	0	0	1	1
slottet	castle	0	0	1	0
slottet	the castle	0	0	1	0
finger	finger	0	0	1	1
finger	finder	0	0	1	0
allra	very	0	0	1	1
allra	most	0	0	1	0
allra	-most; most	0	0	1	0
mun	oral	0	0	1	0
mun	mouth	0	0	1	1
herding	herding	0	0	1	0
seder	seder	0	0	1	0
seder	subsequently	0	0	1	0
seder	custom	0	0	1	0
betonar	stress	0	0	1	0
betonar	emphasize	0	0	1	0
nämnda	said	0	0	1	0
maniska	manic	0	0	1	0
maniska	maniac	0	0	1	0
seden	the seed	0	0	1	0
seden	custom	0	0	1	0
utgåvor	editions	0	0	1	0
utgåvor	issues	0	0	1	0
bildriksdagsval	image election	0	0	1	0
länderna	states	0	0	1	0
länderna	the countries	0	0	1	0
nummer	number	0	0	1	1
store	great	0	0	1	0
kreativitet	creativity	0	0	1	1
autonomi	autonomy	0	0	1	1
trött	tired	0	0	1	1
anfall	attack	0	0	1	1
verka	seem	0	0	1	1
verka	operate	0	0	1	0
verka	appear	0	0	1	1
misshandel	assault	0	0	1	0
misshandel	abuse	0	0	1	0
avrättning	execution	0	0	1	1
farliga	dangerous	0	0	1	0
förslag	proposal	0	0	1	1
förslag	'proposal	0	0	1	0
förslag	proposed	0	0	1	0
allierades	allied's	0	0	1	0
allierades	allied	0	0	1	0
mätningar	measurements	0	0	1	0
mätningar	measurments	0	0	1	0
viruset	virus	0	0	1	0
katarina	katarina	0	0	1	0
hitler	hitler	0	0	1	0
ställning	position	0	0	1	1
ställning	stall	0	0	1	0
solljus	sun light	0	0	1	0
solljus	sunlight	0	0	1	1
skapades	generated	0	0	1	0
skapades	created	0	0	1	0
grundaren	the founder	0	0	1	0
grundaren	founder	0	0	1	0
julian	julian	0	0	1	0
hastighet	speed	0	0	1	1
valt	chosen	0	0	1	0
valt	selected	0	0	1	0
homosexuell	homosexual	0	0	1	1
skalan	scale	0	0	1	0
à	à	0	0	1	0
à	river	0	0	1	0
modernare	mor modern	0	0	1	0
modernare	more modern	0	0	1	0
spritt	spread	0	0	1	0
turistmål	tourist destination	0	0	1	0
turistmål	tourist attraction	0	0	1	0
alltjämt	remains	0	0	1	0
älskade	loved	0	0	1	0
älskade	loved; beloved	0	0	1	0
invasionen	invasion	0	0	1	0
invasionen	the invasion	0	0	1	0
dödad	killed	0	0	1	0
traditionella	traditional	0	0	1	0
traditionella	conventional	0	0	1	0
medlem	member	0	0	1	1
försvinna	vanish	0	0	1	1
försvinna	disappear	0	0	1	1
n	n	0	0	1	0
petrus	petrus	0	0	1	0
schizofreni	schizophrenia	0	0	1	1
depp	depp	0	0	1	0
claes	claes	0	0	1	0
fästning	fastening	0	0	1	0
fästning	fortress	0	0	1	1
della	della	0	0	1	0
nationer	nations	0	0	1	0
tillfällig	temporarily	0	0	1	0
darwins	darwin	0	0	1	0
darwins	darwins	0	0	1	0
vojvodskap	voivodships	0	0	1	0
vojvodskap	voivodeship	0	0	1	0
återvända	return	0	0	1	1
brott	breach	0	0	1	1
brott	crimes	0	0	1	0
brott	crime	0	0	1	1
nationen	the nation	0	0	1	0
kartan	the map	0	0	1	0
kartan	map	0	0	1	0
varefter	whereafter	0	0	1	0
ekonomin	the economy	0	0	1	0
ekonomin	economy	0	0	1	0
traditionellt	traditional	0	0	1	0
ernman	ernman	0	0	1	0
pekar	points	0	0	1	0
pekar	pointer	0	0	1	0
pekar	pointing	0	0	1	0
stadigt	steadily	0	0	1	0
stadigt	stable	0	0	1	0
ersatte	substituting	0	0	1	0
ersatte	replaced	0	0	1	0
pekat	pointed	0	0	1	0
pekat	identified	0	0	1	0
negativ	negative	0	0	1	1
welsh	welsh	0	0	1	0
hundra	hundred	0	0	1	1
hundra	one hundred	0	0	1	0
ändamål	object	0	0	1	1
ändamål	purpose	0	0	1	1
formatet	the format	0	0	1	0
formatet	format	0	0	1	0
formatet	size	0	0	1	0
ersatts	replaced	0	0	1	0
ersatts	(has been) replaced	0	0	1	0
generalguvernören	governor-general	0	0	1	0
generalguvernören	governor general	0	0	1	0
generalguvernören	general governor	0	0	1	0
yngsta	youngest	0	0	1	0
yngste	youngest	0	0	1	0
uppsving	boost	0	0	1	0
gudom	deity	0	0	1	1
dylan	dylan	0	0	1	0
generna	genes	0	0	1	0
generna	the genes	0	0	1	0
charlie	charlie	0	0	1	0
spelad	played	0	0	1	0
handelsmän	merchants	0	0	1	0
förändrats	changed	0	0	1	0
svavel	sulfur	0	0	1	1
svavel	sulphur	0	0	1	1
kemikalier	chemicals	0	0	1	1
fattigare	poorer	0	0	1	0
västsahara	western sahara	0	0	1	0
jean	jean	0	0	1	0
motsatt	opposite	0	0	1	1
motsats	contrary	0	0	1	1
spelar	column	0	0	1	0
spelar	gaming	0	0	1	0
tänkte	thought	0	0	1	0
tänkte	was going to	0	0	1	0
mytologin	mythology	0	0	1	0
kraftigt	heavily	0	0	1	1
torah	torah	0	0	1	1
graden	rate	0	0	1	0
graden	the degree	0	0	1	0
graden	degree	0	0	1	0
europaparlamentet	european-parliament	0	0	1	0
europaparlamentet	the european parliament	0	0	1	0
europaparlamentet	european parliament	0	0	1	0
grader	degrees	0	0	1	0
engelskans	english	0	0	1	0
lärjungar	disciple	0	0	1	0
lärjungar	disciples	0	0	1	0
juridiska	juridical	0	0	1	0
juridiska	legal	0	0	1	0
kalifornien	california	0	0	1	1
gavs	was	0	0	1	0
gavs	gave	0	0	1	0
dödar	kill	0	0	1	0
dödar	kills	0	0	1	0
dödas	put to death	0	0	1	0
dödas	killed	0	0	1	0
dödat	killed	0	0	1	0
eld	fire	0	0	1	1
befälhavare	commander	0	0	1	1
reglera	controlling	0	0	1	0
reglera	expell	0	0	1	0
aktiv	active	1	1	1	1
umeå	umeå	0	0	1	0
regionerna	regions	0	0	1	0
råder	advises	0	0	1	0
råder	is	0	0	1	0
råder	(that) prevails	0	0	1	0
sällskap	company	0	0	1	1
sällskap	groups	0	0	1	0
länk	link	0	0	1	1
enlighet	union	0	0	1	1
enlighet	according (to)	0	0	1	0
enlighet	according	0	0	1	0
rådet	the council	0	0	1	0
rådet	council	0	0	1	0
nobelpriset	the nobel prize	0	0	1	0
nobelpriset	nobel award	0	0	1	0
väljer	elects	0	0	1	0
väljer	select	0	0	1	0
donau	donau	0	0	1	0
donau	danube	0	0	1	0
donau	the danube	0	0	1	0
protesterade	protested	0	0	1	0
auktoritet	authority	0	0	1	1
öronen	lugs	0	0	1	0
öronen	the ears	0	0	1	0
läns	county	0	0	1	0
läns	county's	0	0	1	0
gift	married	0	0	1	1
ladda	load	0	0	1	1
kazakstan	kazakstan	0	0	1	0
kazakstan	kazakhstan	0	0	1	0
ifrån	off	0	0	1	0
bosnienhercegovina	bosnia-hercegovina	0	0	1	0
specifik	specific	0	0	1	1
fotbollen	soccer	0	0	1	0
fotbollen	football	0	0	1	0
hund	dog	0	0	1	1
gifter	marries	0	0	1	0
gifter	toxins	0	0	1	0
lagstiftningen	law-making	0	0	1	0
lagstiftningen	legislation	0	0	1	0
sjöarna	the lakes	0	0	1	0
sjöarna	lakes	0	0	1	0
även	even	0	0	1	1
även	also	0	0	1	1
varianterna	variants	0	0	1	0
varianterna	the diversities	0	0	1	0
hanhon	he/she	0	0	1	0
hanhon	male-female	0	0	1	0
jennifer	jennifer	0	0	1	0
malaysia	malaysia	0	0	1	1
donald	donald	0	0	1	0
xbox	xbox	0	0	1	0
finna	found	0	0	1	0
motsatsen	the opposite	0	0	1	0
motsatsen	opposite	0	0	1	0
vår	spring	0	0	1	1
vår	was	0	0	1	0
området	the area	0	0	1	0
området	area	0	0	1	0
totalt	total	0	0	1	0
totalt	complete	0	0	1	0
totalt	wholly	0	0	1	0
icd	icd	0	0	1	0
våg	vague	0	0	1	0
våg	road	0	0	1	0
våg	wave	0	0	1	1
diktatur	dictator	0	0	1	0
diktatur	dictatorship	0	0	1	1
utse	appoint	0	0	1	0
utse	name	0	0	1	1
enade	united	0	0	1	0
totala	total	0	0	1	0
områden	area	0	0	1	0
områden	areas	0	0	1	0
värd	vard	0	0	1	0
värd	host	0	0	1	1
värd	worth	0	0	1	1
elitserien	elite series	0	0	1	0
elitserien	elitserien	0	0	1	0
uppstått	arised	0	0	1	0
uppstått	resulting	0	0	1	0
uppstått	arisen	0	0	1	0
monoteism	monotheism	0	0	1	1
ishockeyspelare	hockey player	0	0	1	0
ishockeyspelare	ice hockey player	0	0	1	1
ishockeyspelare	hockey players	0	0	1	0
galleri	gallery	0	0	1	1
värt	worth	0	0	1	0
tillbringar	spends	0	0	1	0
tillbringar	spend	0	0	1	0
spelare	player	0	0	1	1
hotellet	the hotel	0	0	1	0
hotellet	hotel	0	0	1	0
meyer	meyer	0	0	1	0
census	census	0	0	1	1
titeln	the title	0	0	1	0
titeln	title	0	0	1	0
tvingades	forced	0	0	1	0
tvingades	had	0	0	1	0
systrar	sisters	0	0	1	0
frälsning	salvation	0	0	1	1
rättvisa	justice	0	0	1	1
plus	plus	0	0	1	1
internationell	international	0	0	1	1
tydliga	clear	0	0	1	0
tydliga	obvious	0	0	1	0
primitiva	primitive	0	0	1	0
civil	civil	0	0	1	1
civil	civilian	0	0	1	1
mörk	dark	0	0	1	1
menade	meant	0	0	1	0
menade	said	0	0	1	0
systemet	the system	0	0	1	0
systemet	system	0	0	1	0
tydligt	clear	0	0	1	0
tydligt	obvious	0	0	1	0
isberg	ice berg	0	0	1	0
isberg	iceberg	0	0	1	1
sinne	mind	0	0	1	1
anorexia	anorexia	0	0	1	0
omges	surrounded	0	0	1	0
omger	surrounds	0	0	1	0
omger	surrounding	0	0	1	0
omger	surrounding the	0	0	1	0
lagt	laid	0	0	1	0
lagt	added	0	0	1	0
kjell	kjell	0	0	1	0
nå	access	0	0	1	0
nå	reach	0	0	1	1
sicilien	sicily	0	0	1	1
västbanken	the west bank	0	0	1	0
västbanken	westbank	0	0	1	0
kronprinsessan	crown princess	0	0	1	0
förtjust	fond	0	0	1	0
förtjust	delighted	0	0	1	1
arbetslösheten	unemployment	0	0	1	0
världsrekord	world record	0	0	1	1
metabolism	metabolism	0	0	1	0
wittenberg	wittenberg	0	0	1	0
dialekterna	dialects	0	0	1	0
fadern	the father	0	0	1	0
skulden	the debt	0	0	1	0
skulden	the guilt	0	0	1	0
italien	italy	0	0	1	1
kingston	kingston	0	0	1	0
människans	humans	0	0	1	0
människans	mankinds	0	0	1	0
människans	human	0	0	1	0
isolering	isolation	0	0	1	1
finns	is	0	0	1	0
finns	exist	0	0	1	0
finns	there is	0	0	1	0
världskrigen	the world wars	0	0	1	0
världskrigen	world wars	0	0	1	0
löser	solve	0	0	1	0
löser	solves	0	0	1	0
eventuell	any	0	0	1	1
fusionen	merger	0	0	1	0
fusionen	the fusion	0	0	1	0
förstå	understandable	0	0	1	0
förstå	understand	0	0	1	1
förstå	first	0	0	1	0
amerikanerna	americans	0	0	1	0
amerikanerna	the americans	0	0	1	0
ruiner	ruins	0	0	1	0
hänga	hang	0	0	1	1
tillika	also	0	0	1	0
tillika	well	0	0	1	0
araber	arabs	0	0	1	0
varifrån	from where; wherefrom	0	0	1	0
varifrån	from which	0	0	1	0
trio	trio	0	0	1	1
bildt	bildt	0	0	1	0
bröstet	chest; breast	0	0	1	0
bröstet	breast	0	0	1	0
döpt	named	0	0	1	0
döpt	baptized	0	0	1	0
öppen	open	0	0	1	1
everest	everest	0	0	1	0
höjer	rises	0	0	1	0
höjer	raise	0	0	1	0
höjer	raising	0	0	1	0
öppet	open	0	0	1	0
hamn	harbor	0	0	1	1
hamn	port	0	0	1	1
hamn	harbour	0	0	1	1
tronen	throne	0	0	1	0
tronen	the throne	0	0	1	0
kambodja	cambodians	0	0	1	0
liberalism	liberalism	0	0	1	1
ni	you	0	0	1	1
margareta	margareta	0	0	1	0
no	no.	0	0	1	0
tillverkade	manufactured	0	0	1	0
tillverkade	made	0	0	1	0
when	when	0	0	1	0
nf	nf	0	0	1	0
saturnus	saturn	0	0	1	1
saturnus	saturnus	0	0	1	0
läkemedel	drugs	0	0	1	0
läkemedel	medicine	0	0	1	1
ny	new	0	0	1	1
tio	ten	0	0	1	1
tid	time	0	0	1	1
nr	no.	0	0	1	0
nr	number	0	0	1	0
nr	no	0	0	1	0
nivå	niva	0	0	1	0
nivå	level	0	0	1	1
nu	now	0	0	1	1
picture	picture	0	0	1	0
phoenix	phoenix	0	0	1	0
erhållit	obtained	0	0	1	0
erhållit	acquired	0	0	1	0
erhållit	received	0	0	1	0
källkod	source	0	0	1	0
källkod	source code	0	0	1	0
football	football	0	0	1	0
miscellaneous	miscellaneous	0	0	1	0
romersk	roman	0	0	1	1
tunna	thin	0	0	1	0
massakern	massacre	0	0	1	0
estetik	stetik	0	0	1	0
estetik	esthetics	0	0	1	0
estetik	aesthetics	0	0	1	1
förväxlas	mistaken	0	0	1	0
förväxlas	confused	0	0	1	0
förväxlas	mixed up (with)	0	0	1	0
utrustning	equipment	0	0	1	1
utrustning	gear	0	0	1	0
ultraviolett	ultraviolet	0	0	1	1
ovanstående	above	0	0	1	1
ovanstående	previously instructed	0	0	1	0
lördagen	the saturday	0	0	1	0
lördagen	saturday	0	0	1	0
första	first	0	0	1	1
förste	chief	0	0	1	1
förste	the first	0	0	1	0
förste	first	0	0	1	1
beroendeframkallande	addictive	0	0	1	0
vietnam	vietnam	0	0	1	1
cellens	the cell's	0	0	1	0
cellens	cell's	0	0	1	0
cellens	the cells	0	0	1	0
påbörjade	started	0	0	1	0
påbörjade	began	0	0	1	0
rom	rome	0	0	1	1
rom	rom	0	0	1	0
ron	ron	0	0	1	0
rob	rob	0	0	1	0
fördelar	share	0	0	1	0
fördelar	advantages	0	0	1	0
fördelar	advantage	0	0	1	0
övergripande	over arching	0	0	1	0
övergripande	overall	0	0	1	0
övergripande	general	0	0	1	0
josé	jose	0	0	1	0
roy	roy	0	0	1	0
koreanska	korean	0	0	1	0
tillgänglig	available	0	0	1	1
tillgänglig	provided	0	0	1	0
udda	odd	0	0	1	1
minska	reducing	0	0	1	0
minska	reduce	0	0	1	1
förändrades	changed	0	0	1	0
hundraser	breeds	0	0	1	0
hundraser	alternative strains	0	0	1	0
hundraser	breed of dogs	0	0	1	0
laura	laura	0	0	1	0
kallar	call	0	0	1	0
kallar	calls	0	0	1	0
mottagarens	the reciever	0	0	1	0
mottagarens	the receivers	0	0	1	0
mottagarens	the receiver's	0	0	1	0
bägge	both	0	0	1	0
bägge	ram	0	0	1	0
ständerna	the cities	0	0	1	0
konstitutionell	constitutional	0	0	1	1
tanke	light	0	0	1	0
tanke	in light of	0	0	1	0
federation	federation	0	0	1	1
försvarsminister	minister of defence	0	0	1	0
varvid	in which	0	0	1	0
flytt	escaped	0	0	1	0
flytt	move	0	0	1	0
flytt	fled	0	0	1	0
krossa	crush	0	0	1	1
krossa	crushing	0	0	1	0
metod	method	0	0	1	1
hawaii	hawaii	0	0	1	0
begränsa	limit	0	0	1	1
christmas	christmas	0	0	1	0
olyckor	accidents	0	0	1	0
lever	living	0	0	1	0
lever	live	0	0	1	0
lever	liver	0	0	1	1
der	where	0	0	1	0
der	german word	0	0	1	0
höga	high	0	0	1	0
heinz	heinz	0	0	1	0
trend	trend	0	0	1	1
stilar	styles	0	0	1	0
kategorirock	category:rock	0	0	1	0
kategorirock	category rock	0	0	1	0
colin	colin	0	0	1	0
högt	high	0	0	1	1
högt	highly	0	0	1	0
port	gate	0	0	1	1
port	port	0	0	1	0
uppgifterna	data	0	0	1	0
uppgifterna	the information	0	0	1	0
tillhörde	was a part of	0	0	1	0
tillhörde	belonging to	0	0	1	0
tillhörde	belonged to	0	0	1	0
bilmärke	car make	0	0	1	0
bilmärke	make of car	0	0	1	0
bestå	consists	0	0	1	0
bestå	exist	0	0	1	0
bestå	comprise	0	0	1	0
poesi	poetry	0	0	1	1
övertalade	over spoke	0	0	1	0
övertalade	persuaded	0	0	1	0
miniatyr	miniature	0	0	1	1
miniatyr	thumbnail	0	0	1	0
ingenjör	engineering	1	1	0	0
ingenjör	complex	1	0	1	0
ingenjör	hard	1	0	1	0
ingenjör	ingenjor	1	0	1	0
ingenjör	engineer	1	1	0	1
åtgärder	measures	0	0	1	0
angelina	angelina	0	0	1	0
gravitation	gravitation	0	0	1	1
gravitation	gravity	0	0	1	1
kamp	struggle	0	0	1	1
kamp	fight	0	0	1	1
vindkraftverk	wind turbine	0	0	1	0
vindkraftverk	wind power station	0	0	1	0
enkla	simple	0	0	1	0
enkla	single	0	0	1	0
premiärminister	prime minister	0	0	1	1
metaller	metals	0	0	1	0
utåt	outwardly	0	0	1	1
utåt	out	0	0	1	0
jord	soil	0	0	1	1
jord	earth	0	0	1	1
turister	tourists	0	0	1	0
dublin	dublin	0	0	1	0
lokal	local	0	0	1	1
ankomst	arrival	0	0	1	1
experimenterade	experimented	0	0	1	0
tilltagande	increasing	0	0	1	1
barndom	childhood	0	0	1	1
rafael	rafael	0	0	1	0
rafael	rafel	0	0	1	0
framför	in front of	0	0	1	1
framför	particularly	0	0	1	0
framför	above	0	0	1	1
luften	air	0	0	1	0
sikt	term	0	0	1	1
sikt	run	0	0	1	1
sikt	sit	0	0	1	0
tillfälliga	temporary	0	0	1	0
etablera	erablera	0	0	1	0
etablera	establish	0	0	1	1
etablera	up	0	0	1	0
trummor	drums	0	0	1	0
tillfälligt	temporarly	0	0	1	0
tillfälligt	temporary	0	0	1	0
bolaget	company	0	0	1	0
bolaget	the company	0	0	1	0
ungerska	hungarian	0	0	1	1
härskare	ruler	0	0	1	1
undan	away (from)	0	0	1	0
undan	escape	0	0	1	0
utropades	proclaimed	0	0	1	0
utropades	was proclaimed	0	0	1	0
samfundet	the communion	0	0	1	0
samfundet	association	0	0	1	0
begå	commit	0	0	1	1
anda	spirit	0	0	1	1
begäran	request	0	0	1	1
inblandade	involved	0	0	1	0
andy	andy	0	0	1	0
kurder	kurds	0	0	1	0
australian	australian	0	0	1	0
utgåvan	edition	0	0	1	0
utgåvan	the edition	0	0	1	0
utgåvan	issue	0	0	1	0
uppskattningar	estimates	0	0	1	0
typerna	the types	0	0	1	0
typerna	types	0	0	1	0
författningen	constitution	0	0	1	0
palestinsk	palestinian	0	0	1	1
inbördeskrig	civil war	0	0	1	1
efterhand	post	0	0	1	0
efterhand	hindsight	0	0	1	0
piano	piano	0	0	1	1
styras	guided	0	0	1	0
styras	controlled	0	0	1	0
styras	steered	0	0	1	0
drabbades	affected	0	0	1	0
drabbades	where hit by	0	0	1	0
drabbades	afflicted	0	0	1	0
julius	julius	0	0	1	0
musikaliska	musical	0	0	1	0
valla	herd	0	0	1	1
valla	valla	0	0	1	0
valla	wax	0	0	1	0
jude	dude	0	0	1	0
jude	jew	0	0	1	1
allvarlig	serious	0	0	1	1
judy	judy	0	0	1	1
humle	hops	0	0	1	0
humle	hop	0	0	1	1
generell	general	0	0	1	1
befolkningstäthet	population density	0	0	1	1
befolkningstäthet	the population density	0	0	1	0
karibiska	caribbean	0	0	1	0
musikaliskt	musically talented	0	0	1	0
musikaliskt	musical	0	0	1	0
musikaliskt	musically	0	0	1	0
springsteens	springsteen's	0	0	1	0
springsteens	springsteens	0	0	1	0
dokumenterade	documented	0	0	1	0
utdelades	distributed	0	0	1	0
utdelades	awarded	0	0	1	0
hemligt	secret	0	0	1	0
annorlunda	different	0	0	1	0
annorlunda	otherwise	0	0	1	1
hemliga	secret	0	0	1	0
swedish	swedish	0	0	1	0
omvända	reverse	0	0	1	0
hört	heard	0	0	1	0
hört	heared	0	0	1	0
frivilligt	voluntarily	0	0	1	0
frivilligt	voluntary	0	0	1	0
sydöst	south east	0	0	1	0
sydöst	southeast	0	0	1	1
frivilliga	volunteers	0	0	1	0
frivilliga	optional	0	0	1	0
frivilliga	voluntary	0	0	1	0
andlig	spiritual	0	0	1	1
andlig	spirtual	0	0	1	0
simning	swimming	0	0	1	1
regeln	the rule	0	0	1	0
regeln	rule	0	0	1	0
muslimerna	muslims	0	0	1	0
muslimerna	the muslims	0	0	1	0
inriktad	focused on	0	0	1	0
inriktad	oriented	0	0	1	0
inriktad	intent	0	0	1	0
etablerat	established	0	0	1	0
tillfälle	instance	0	0	1	0
tillfälle	occasion	0	0	1	1
tillfälle	time	0	0	1	0
tvserien	tv series	0	0	1	0
tvserien	the tv show	0	0	1	0
tvserien	television program	0	0	1	0
levt	survived	0	0	1	0
fascism	fascism	0	0	1	1
sydliga	southern	0	0	1	0
tvserier	tv-shows	0	0	1	0
tvserier	tv shows	0	0	1	0
tvserier	tv-series	0	0	1	0
belagt	coated	0	0	1	0
fenomen	phenomena	0	0	1	0
fenomen	phenomenon	0	0	1	1
fenomen	phenomenazaqq	0	0	1	0
leva	live	0	0	1	1
utrikespolitiska	foreign policy	0	0	1	0
utrikespolitiska	foreign political	0	0	1	0
berättar	tells	0	0	1	0
berättas	(as) told	0	0	1	0
berättas	is told	0	0	1	0
berättas	told	0	0	1	0
berättat	told	0	0	1	1
marknad	market	0	0	1	1
kroniska	chronic	0	0	1	0
beror	is	0	0	1	0
stridande	fighting	0	0	1	1
stridande	conflict	0	0	1	0
stridande	warring	0	0	1	0
japanska	japanese	0	0	1	0
anlände	arrived	0	0	1	0
förknippas	associated to	0	0	1	0
förknippas	associated	0	0	1	0
förknippas	associate	0	0	1	0
representation	representation	0	0	1	1
kategoriamerikanska	u.s. category	0	0	1	0
pappa	dad	0	0	1	1
komplicerad	complex	0	0	1	1
komplicerad	complicated	0	0	1	1
följden	the result	0	0	1	0
följden	the cause	0	0	1	0
följden	result	0	0	1	0
idéerna	ideema	0	0	1	0
idéerna	ideas	0	0	1	0
orter	varieties	0	0	1	0
orter	locations	0	0	1	0
kartor	maps	0	0	1	0
bushs	bush's	0	0	1	0
bushs	bush	0	0	1	0
orten	resort	0	0	1	0
orten	the suburb	0	0	1	0
släktet	the genus	0	0	1	0
följder	impact	0	0	1	0
följder	consequences	0	0	1	0
behövs	required	0	0	1	0
behövs	is needed	0	0	1	0
komplicerat	complex	0	0	1	0
komplicerat	complicated	0	0	1	0
iberiska	iberian	0	0	1	0
fasen	phase	0	0	1	0
rapport	report	0	0	1	1
wallace	wallace	0	0	1	0
utvecklingen	development	0	0	1	0
utvecklingen	the development	0	0	1	0
organisation	body	0	0	1	0
organisation	organization	0	0	1	1
sträcker	stretches	0	0	1	0
sträcker	extend	0	0	1	0
behandlingen	the treatment	0	0	1	0
behandlingen	the treament	0	0	1	0
behandlingen	treatment	0	0	1	0
energikälla	source	0	0	1	0
energikälla	energy source	0	0	1	0
energikälla	energy call	0	0	1	0
spelarna	players	0	0	1	0
klassen	the class	0	0	1	0
klassen	klasses	0	0	1	0
pågående	current	0	0	1	0
pågående	ongoing	0	0	1	1
marleys	marley's	0	0	1	0
marleys	marley	0	0	1	0
passar	suitable	0	0	1	0
passar	suits	0	0	1	0
femte	fifth	0	0	1	1
övertyga	convince	0	0	1	1
övertyga	convince our	0	0	1	0
hamilton	hamilton	0	0	1	0
karlsson	karlsson	0	0	1	0
tredjedel	tredjedel	0	0	1	0
tredjedel	a third	0	0	1	0
tredjedel	third	0	0	1	1
hotar	threatens	0	0	1	0
term	term	0	0	1	1
dåligt	poor	0	0	1	0
opera	opera	0	0	1	1
opera	operator	0	0	1	0
ägda	owned	0	0	1	0
snabb	instant	0	0	1	0
ägde	tookplace; occured	0	0	1	0
ägde	was	0	0	1	0
ägde	owned	0	0	1	0
futharkens	futharkens	0	0	1	0
futharkens	futhark	0	0	1	0
futharkens	the futhark's	0	0	1	0
viggo	viggo	0	0	1	0
alternativ	alternative	0	0	1	1
hotad	threatened	0	0	1	0
nöjd	content	0	0	1	1
bildning	education	0	0	1	1
bildning	form	0	0	1	1
bildning	learning	0	0	1	1
semifinal	semifinals	0	0	1	0
semifinal	semi finals	0	0	1	0
stressorer	stressors	0	0	1	0
dömd	sentenced	0	0	1	0
dömd	convicted	0	0	1	0
hoppade	jumped	0	0	1	0
tänka	thinking	0	0	1	0
tänka	think	0	0	1	1
tänka	fill	0	0	1	0
besöker	visit	0	0	1	0
besöker	visits	0	0	1	0
läggas	laid	0	0	1	0
läggas	added	0	0	1	0
tänkt	expected	0	0	1	0
tänkt	supposed; intended	0	0	1	0
tänkt	intended	0	0	1	0
amerikansk	american	0	0	1	1
amerikansk	u.s.	0	0	1	0
behandlar	treats	0	0	1	0
behandlar	treat	0	0	1	0
behandlas	treated	0	0	1	0
upprepade	repeated	0	0	1	0
accepterad	acceptable	0	0	1	0
stortorget	stortorget	0	0	1	0
stortorget	the main square	0	0	1	0
profil	profile	0	0	1	1
accepterar	accepts	0	0	1	0
accepterar	accept	0	0	1	0
accepterat	accepted	0	0	1	0
kent	kent	0	0	1	0
utlösa	trigger	0	0	1	0
brett	broad	0	0	1	0
juldagen	christmas day	0	0	1	1
zuckerberg	zuckerberg	0	0	1	0
etanol	ethanol	0	0	1	1
hjalmar	hjalmar	0	0	1	0
gallien	gaul	0	0	1	1
avtalet	the treaty	0	0	1	0
avtalet	the contract	0	0	1	0
avtalet	agreement	0	0	1	0
arbetet	work	0	0	1	0
arbetet	the work	0	0	1	0
traditionen	the tradition	0	0	1	0
traditionen	tradition	0	0	1	0
motion	motion	0	0	1	1
motion	exercise	0	0	1	1
traditioner	traditions	0	0	1	0
traditioner	the traditions	0	0	1	0
place	place	0	0	1	0
politiken	policy	0	0	1	0
politiken	the politics	0	0	1	0
hemsida	website	0	0	1	0
hemsida	homepage	0	0	1	0
blood	blood	0	0	1	0
origin	origin	0	0	1	0
rené	rené	0	0	1	0
rené	rene	0	0	1	0
george	george	0	0	1	0
respekt	respected	0	0	1	0
respekt	respect	0	0	1	1
given	given	0	0	1	1
ian	ian	0	0	1	0
skjuten	shot	0	0	1	0
anderson	anderson	0	0	1	0
bahamas	bahamas	0	0	1	0
österrikes	austria's	0	0	1	0
österrikes	austrias	0	0	1	0
skjuter	shoots	0	0	1	0
skjuter	slide	0	0	1	0
skjuter	extend	0	0	1	0
givet	granted	0	0	1	0
givet	given	0	0	1	0
hud	skin	0	0	1	1
spelats	been played	0	0	1	0
spelats	recorded	0	0	1	0
spelats	played	0	0	1	0
webbplatser	webbsites	0	0	1	0
webbplatser	websites	0	0	1	0
gia	gia	0	0	1	0
grund	because	0	0	1	0
grund	in the context: "på grund" = because of	0	0	1	0
montenegro	montenergo	0	0	1	0
montenegro	montenegro	0	0	1	0
alan	alan	0	0	1	0
kallade	called	0	0	1	0
håkan	chin	0	0	1	0
håkan	håkan	0	0	1	0
hur	how	0	0	1	1
hur	the	0	0	1	0
hur	cage	0	0	1	0
hus	house	0	0	1	1
hus	housing	0	0	1	1
hus	a house	0	0	1	0
webbplatsen	webpage	0	0	1	0
webbplatsen	the website	0	0	1	0
webbplatsen	site	0	0	1	0
population	population	0	0	1	0
smeknamn	nickname	0	0	1	0
officerare	officers	0	0	1	0
officerare	officer	0	0	1	0
modellen	model	0	0	1	0
modellen	the model	0	0	1	0
balans	balance	0	0	1	1
marinen	navy	0	0	1	0
marinen	marines	0	0	1	0
kontroll	control	0	0	1	1
spänning	voltage	0	0	1	1
r	r	0	0	1	0
modeller	models	0	0	1	0
beräknar	calculates the	0	0	1	0
beräknar	computes	0	0	1	0
beräknar	values	0	0	1	0
bildades	founded	0	0	1	0
bildades	formed	0	0	1	0
bildades	was formed	0	0	1	0
rena	pure	0	0	1	0
mottagare	recipient	0	0	1	1
mottagare	receiver	0	0	1	1
nätvingar	it's a animal	1	0	1	0
nätvingar	natvinger	1	0	1	0
nätvingar	net wings	1	0	1	0
nätvingar	lacewings	1	0	1	0
nätvingar	each	1	0	1	0
nätvingar	net-winged insects	1	1	0	0
nätvingar	night wings	1	1	0	0
nätvingar	neuropteran	1	0	1	0
nätvingar	neuropterans	1	1	0	0
nätvingar	neuroptera	1	1	0	0
nätvingar	(nätvingar) an order in the class insects.	1	0	1	0
nätvingar	nätvingar	1	0	1	0
nätvingar	netwings	1	0	1	0
nätvingar	lacewing	1	0	1	0
nätvingar	natvingar	1	0	1	0
ana	feel	0	0	1	0
ana	ana	0	0	1	0
lösningen	the solution	0	0	1	0
lösningen	solution	0	0	1	0
hållit	held	0	0	1	0
hållit	maintained	0	0	1	0
hållit	kept	0	0	1	0
kromosomerna	chromosomes	0	0	1	0
kromosomerna	the chromosomes	0	0	1	0
maten	the food	0	0	1	0
mando	command	0	0	1	0
rent	true	0	0	1	0
rent	clean	0	0	1	0
jordskorpan	earth's crust	0	0	1	0
jordskorpan	earth crust	0	0	1	0
jordskorpan	the earth's crust	0	0	1	0
malta	malta	0	0	1	1
ideal	ideals	0	0	1	0
ideal	ideal	0	0	1	1
gustavs	gustavs	0	0	1	0
gustavs	gustav	0	0	1	0
konsert	concert	0	0	1	1
periodvis	periodically	0	0	1	0
vårt	our	0	0	1	0
vårt	each	0	0	1	0
knutna	attached	0	0	1	0
knutna	associated	0	0	1	0
knutna	tied	0	0	1	0
våra	our	0	0	1	0
släktingar	relatives	0	0	1	0
målvakt	goalee	0	0	1	0
målvakt	goalkeeper	0	0	1	1
vård	vard	0	0	1	0
vård	nursing	0	0	1	0
vård	healthcare	0	0	1	0
diskussioner	discussions	0	0	1	0
diskussioner	discussion	0	0	1	0
biogeografi	biogeography	1	1	0	0
biogeografi	evolution	1	0	1	0
biogeografi	use	1	0	1	0
biogeografi	biogegraphy	1	0	1	0
biogeografi	usage	1	0	1	0
biogeografi	biogeografi	1	0	1	0
falla	fall	0	0	1	1
fria	free	0	0	1	0
ledamöter	commissioners	0	0	1	0
ledamöter	members	0	0	1	0
staterna	states	0	0	1	0
staterna	usa	0	0	1	0
lisbet	lisbet	0	0	1	0
astronomiska	astronomical	0	0	1	0
betydande	important	0	0	1	1
betydande	significant	0	0	1	0
utkämpades	fought	0	0	1	0
herren	lord	0	0	1	0
herren	the lord	0	0	1	1
målet	minced	0	0	1	0
målet	target	0	0	1	0
målet	the target	0	0	1	0
frågan	issue	0	0	1	0
frågan	the question	0	0	1	0
tron	faith	0	0	1	0
djur	animals	0	0	1	0
djur	animal	0	0	1	1
ronaldinho	ronaldinho	0	0	1	0
förlopp	process	0	0	1	0
förlopp	pattern	0	0	1	1
förlopp	developments	0	0	1	0
framgångarna	successes	0	0	1	0
framgångarna	the successes	0	0	1	0
sjunka	decrease	0	0	1	0
sjunka	descend	0	0	1	1
tror	believe	0	0	1	0
tror	think	0	0	1	0
bandets	the bands	0	0	1	0
bandets	band	0	0	1	0
räcker	enough	0	0	1	0
räcker	sufficient	0	0	1	0
gula	yellow	0	0	1	0
tvprogram	tv program	0	0	1	0
tvprogram	tv-show	0	0	1	0
guld	gold	0	0	1	1
könen	the sexes	0	0	1	0
könen	equality	0	0	1	0
tidningarna	papers	0	0	1	0
flydde	fled	0	0	1	0
löper	runs	0	0	1	0
löper	at	0	0	1	0
ovanligt	unusual	0	0	1	0
ovanligt	rare	0	0	1	0
gult	yellow	0	0	1	1
matematiska	mathematical	0	0	1	0
ovanliga	unusual	0	0	1	0
ovanliga	rare	0	0	1	0
analys	analysis	0	0	1	1
larsson	larsson	0	0	1	0
aktiviteten	the level of activity	0	0	1	0
aktiviteten	activity	0	0	1	0
grundandet	founding (of)	0	0	1	0
grundandet	founding	0	0	1	0
jazz	jazz	0	0	1	1
administrativ	administration	0	0	1	0
administrativ	administrative	0	0	1	1
forsberg	forsberg	0	0	1	0
tåg	rail	0	0	1	0
tåg	trains	0	0	1	0
beredd	ready (to)	0	0	1	0
beredd	prepared	0	0	1	1
avsåg	meant	0	0	1	0
avsåg	intended	0	0	1	0
avsåg	mean	0	0	1	0
självständig	independent	0	0	1	1
självständig	independently	0	0	1	0
självständig	independant	0	0	1	0
skivkontrakt	record deal	0	0	1	0
skivkontrakt	record contract	0	0	1	0
dramat	drama	0	0	1	0
dramat	the drama	0	0	1	0
joker	joker	0	0	1	1
kommitté	committee	0	0	1	0
republika	republic	0	0	1	0
republika	republika	0	0	1	0
baltikum	the baltics	0	0	1	0
baltikum	baltics	0	0	1	0
satte	put	0	0	1	0
satte	sat	0	0	1	0
satte	put together	0	0	1	0
minnen	memories	0	0	1	0
minnen	memory	0	0	1	0
utsätts	exposed	0	0	1	0
beethoven	beethoven	0	0	1	0
kraftigare	greater	0	0	1	0
kraftigare	more powerfully	0	0	1	0
inspelningen	recording	0	0	1	0
uppdraget	task; assignment	0	0	1	0
uppdraget	assignment	0	0	1	0
finansiering	financing	0	0	1	0
finansiering	financiation	0	0	1	0
tekniskt	technical	0	0	1	0
college	college	0	0	1	1
såldes	sold	0	0	1	0
stanley	stanley	0	0	1	0
minnet	the memory	0	0	1	0
minnet	memory	0	0	1	0
påstod	claimed	0	0	1	0
påstod	said	0	0	1	0
freden	the peace	0	0	1	0
freden	peace	0	0	1	0
federal	federal	0	0	1	1
officiellt	official	0	0	1	0
officiellt	officially	0	0	1	1
utbud	range	0	0	1	0
utbud	availibility	0	0	1	0
utbud	supply	0	0	1	0
skett	done	0	0	1	0
skett	happened	0	0	1	0
därifrån	from thence	0	0	1	1
därifrån	from there	0	0	1	1
för	of	0	0	1	1
för	to; for	0	0	1	0
för	for	0	0	1	1
intresserad	interested	0	0	1	1
mellan	between	0	0	1	1
antagligen	ligands presumably	0	0	1	0
antagligen	probably	0	0	1	1
antagligen	presumably	0	0	1	1
myter	myths	0	0	1	0
ersättare	alternate	0	0	1	0
ersättare	replacement	0	0	1	0
come	come	0	0	1	0
summa	sum	0	0	1	1
summa	total	0	0	1	1
sydeuropa	south europe	0	0	1	0
sydeuropa	southern europe	0	0	1	1
region	region	0	0	1	0
ordagrant	literally	0	0	1	1
ordagrant	literal	0	0	1	0
ordagrant	verbatim	0	0	1	1
spindlar	spiders	0	0	1	0
nöd	distress	0	0	1	1
nöd	emergency	0	0	1	0
diskriminering	discrimination	0	0	1	1
ägare	owner	0	0	1	1
ägare	owners	0	0	1	0
lenins	lenin	0	0	1	0
lenins	lenin's	0	0	1	0
introducerades	introduced	0	0	1	0
gjorde	did	0	0	1	0
gjorda	made	0	0	1	0
gjorda	done	0	0	1	0
pakistan	pakistan	0	0	1	1
behandla	treatment	0	0	1	0
period	period	0	0	1	1
pop	pop	0	0	1	1
försvunnit	disappeared	0	0	1	0
fransk	french	0	0	1	1
fransk	france	0	0	1	0
werner	werner	0	0	1	0
statens	state	0	0	1	0
statens	the government's	0	0	1	0
utformning	formation	0	0	1	1
utformning	shape	0	0	1	1
utformning	layout	0	0	1	0
poe	poe	0	0	1	0
åland	Åland	0	0	1	0
howard	howard	0	0	1	0
folken	the peoples	0	0	1	0
folken	peoples	0	0	1	0
folken	people	0	0	1	0
strikta	strict	0	0	1	0
värde	let there be	0	0	1	0
värde	value	0	0	1	1
stödjer	support	0	0	1	0
stödjer	supports	0	0	1	0
dagarna	the days	0	0	1	0
dagarna	day	0	0	1	0
musikstil	music	0	0	1	0
musikstil	music still	0	0	1	0
musikstil	music style	0	0	1	0
folket	the people	0	0	1	0
folket	people	0	0	1	0
invaderade	invaded	0	0	1	0
anderna	andes	0	0	1	0
anderna	the andes	0	0	1	0
andres	andres	0	0	1	0
andres	other's	0	0	1	0
andrew	andrew	0	0	1	0
kapitulation	surrender	0	0	1	0
kapitulation	capitulation	0	0	1	1
tiger	tiger	0	0	1	1
tiger	silent	0	0	1	0
nivåer	levels	0	0	1	0
minister	minister	0	0	1	1
konstruerade	constructed	0	0	1	0
kaos	chaos	0	0	1	1
andrea	andrea	0	0	1	0
champions	campion	0	0	1	0
champions	champions	0	0	1	0
hughes	hughes	0	0	1	0
odlade	grew	0	0	1	0
odlade	dlade	0	0	1	0
odlade	cultured	0	0	1	0
riktade	targeted	0	0	1	0
bilda	form	0	0	1	1
tillåta	allow to	0	0	1	0
tillåta	allowing	0	0	1	0
tillåta	allow	0	0	1	1
mount	mount	0	0	1	0
influenser	influence	0	0	1	0
influenser	influences	0	0	1	0
cash	cash	0	0	1	0
arnold	arnold	0	0	1	0
spreds	spread	0	0	1	0
spreds	disseminated	0	0	1	0
fiende	enemy	0	0	1	1
föregående	preceeding; previous	0	0	1	0
föregående	previous	0	0	1	1
grundlagen	constitution	0	0	1	0
grundlagen	the constitutional law	0	0	1	0
tillåts	is allowed	0	0	1	0
tillåts	allowed	0	0	1	0
odens	odin's	0	0	1	0
odens	node	0	0	1	0
odens	oden's	0	0	1	0
universums	universe	0	0	1	0
universums	the universe's	0	0	1	0
universums	universe's	0	0	1	0
upprätthålla	maintain	0	0	1	1
upprätthålla	keep up	0	0	1	1
upprätthålla	maintaining	0	0	1	0
sänder	broadcast	0	0	1	0
sänder	transmits	0	0	1	0
sändes	was sent	0	0	1	0
sändes	sent	0	0	1	0
pippi	birdie	0	0	1	0
pippi	pippi	0	0	1	0
knyta	tie	0	0	1	1
gröna	green	0	0	1	0
övertogs	were taken	0	0	1	0
övertogs	overtaken	0	0	1	0
övertogs	over were taken	0	0	1	0
status	status	0	0	1	1
går	is	0	0	1	0
går	goes	0	0	1	0
producera	produce	0	0	1	1
producera	producing	0	0	1	0
republikens	republic's	0	0	1	0
republikens	republic	0	0	1	0
fysiologi	physiology	0	0	1	1
protoner	protons	0	0	1	0
persons	a person's	0	0	1	0
persons	persons	0	0	1	0
persons	person's	0	0	1	0
linjerna	routes	0	0	1	0
linjerna	the lines	0	0	1	0
linjerna	lines	0	0	1	0
köpt	purchased	0	0	1	0
köpt	bought	0	0	1	0
vatikanstaten	vatican city	0	0	1	0
vatikanstaten	the vatican	0	0	1	0
vatikanstaten	vatican	0	0	1	0
relaterade	related	0	0	1	0
mäts	measured	0	0	1	0
mäts	is measured	0	0	1	0
modet	the fashion	0	0	1	0
modet	courage	0	0	1	0
modet	fashion	0	0	1	0
medvetna	conscious	0	0	1	0
medvetna	aware	0	0	1	0
kommunistisk	communistic	0	0	1	1
kommunistisk	communist	0	0	1	1
mätt	measured	0	0	1	1
mätt	dull	0	0	1	0
pennsylvania	pennsylvania	0	0	1	0
breda	broad	0	0	1	0
breda	wide	0	0	1	0
breda	qual o curso que você está estudando	0	0	1	0
mäta	compare	0	0	1	0
mäta	feeding	0	0	1	0
without	without	0	0	1	0
nordkoreas	north korea	0	0	1	0
nordkoreas	north korea's	0	0	1	0
nordkoreas	north coreas	0	0	1	0
kopplingen	the connection	0	0	1	0
kopplingen	coupling	0	0	1	0
lyckan	the happiness	0	0	1	0
lyckan	happiness	0	0	1	0
listorna	menus	0	0	1	0
listorna	the lists of candidates	0	0	1	0
listorna	the lists	0	0	1	0
utländska	foreign	0	0	1	0
övre	upper	0	0	1	1
övre	top	0	0	1	1
kommentarer	comments	0	0	1	0
actress	actress	0	0	1	0
actress	online	0	0	1	0
janukovytj	janukovytj	0	0	1	0
janukovytj	yanukovych	0	0	1	0
ekologiska	ecological	0	0	1	0
enligt	according (to)	0	0	1	0
enligt	according to	0	0	1	1
kill	kill	0	0	1	0
kill	kill found	0	0	1	0
harrison	harrison	0	0	1	0
lyckas	successful	0	0	1	0
lyckas	succeed	0	0	1	1
räkna	count	0	0	1	1
räkna	special	0	0	1	0
leta	search	0	0	1	1
leta	check	0	0	1	0
utvinns	extracted	0	0	1	0
starka	strong	0	0	1	0
tim	tim	0	0	1	0
tim	h	0	0	1	0
rose	rose	0	0	1	0
regent	ruler	0	0	1	0
regent	regent	0	0	1	1
storstäder	metropolises	0	0	1	0
storstäder	cities	0	0	1	0
rosa	pink	0	0	1	1
rosa	rosa	0	0	1	0
utbyte	yield	0	0	1	1
utbyte	trade	0	0	1	1
starkt	strongly	0	0	1	1
starkt	strong	0	0	1	1
lett	resulted	0	0	1	0
lett	led (to)	0	0	1	0
utvinna	extract	0	0	1	1
grupper	groups	0	0	1	0
feminism	feminism	0	0	1	1
ross	ross	0	0	1	0
arméer	armies	0	0	1	0
arméer	army	0	0	1	0
riket	kingdom	0	0	1	0
riket	the land	0	0	1	0
riket	whole country	0	0	1	0
mesta	most	0	0	1	0
vampyren	the vampire	0	0	1	0
vampyren	vampire	0	0	1	0
införandet	introduction	0	0	1	0
införandet	the introduction	0	0	1	0
delhi	delhi	0	0	1	1
utrikespolitik	foreign policy	0	0	1	1
utrikespolitik	foreign affairs	0	0	1	0
utrikespolitik	forgein policy	0	0	1	0
uppslagsordet	lookup word	0	0	1	0
uppslagsordet	lexical entry; word	0	0	1	0
uppslagsordet	entry word	0	0	1	0
kille	guy	0	0	1	1
majoritet	majority	0	0	1	1
inflation	inflation	0	0	1	1
vampyrer	vampires	0	0	1	0
rättigheterna	the rights	0	0	1	0
rättigheterna	rights	0	0	1	0
sådan	such	0	0	1	1
sådan	kind of	0	0	1	0
walk	walk	0	0	1	0
förrän	until	0	0	1	0
förrän	before	0	0	1	1
riken	the kingdoms	0	0	1	0
riken	kingdoms	0	0	1	0
kommentar	comment	0	0	1	1
privilegium	privelege	1	0	1	0
privilegium	oh	1	0	1	0
privilegium	prerogative	1	1	0	1
privilegium	privileium	1	0	1	0
privilegium	privilege	1	1	0	1
privilegium	privlege	1	0	1	0
privilegium	privledge	1	0	1	0
afrikas	africa's	0	0	1	0
afrikas	africas	0	0	1	0
afrikas	africa	0	0	1	0
kennedy	kennedy	0	0	1	0
mexikanska	mexican	0	0	1	0
sverigedemokraterna	sweden democrats	0	0	1	0
sverigedemokraterna	swedish democracy	0	0	1	0
göteborg	gothenburg	0	0	1	1
cooper	cooper	0	0	1	0
tower	tower	0	0	1	0
são	sao	0	0	1	0
rammstein	rammstein	0	0	1	0
tillfället	to the case	0	0	1	0
tillfället	time	0	0	1	0
verksamheten	the work	0	0	1	0
verksamheten	activity	0	0	1	0
madrid	madrid	0	0	1	1
teorin	theory	0	0	1	0
teorin	the theory	0	0	1	0
passera	pass	0	0	1	1
latinet	latin	0	0	1	0
världsarv	world heritage	0	0	1	0
alkoholer	alcohols	0	0	1	0
verksamheter	operations	0	0	1	0
verksamheter	businesses	0	0	1	0
verksamheter	activity	0	0	1	0
tillfällen	jobs	0	0	1	0
tillfällen	occasion	0	0	1	0
tillfällen	oppertunities	0	0	1	0
tiders	days'	0	0	1	0
tiders	time's	0	0	1	0
tiders	times	0	0	1	0
fiktion	fiction	0	0	1	1
inspirerades	(was) inspired	0	0	1	0
inspirerades	inspired	0	0	1	0
sitta	sit	0	0	1	1
stopp	stop	0	0	1	1
moon	moon	0	0	1	0
skära	carve	0	0	1	1
skära	cut	0	0	1	1
skära	army	0	0	1	0
buddha	buddha	0	0	1	1
inträffade	occurred	0	0	1	0
inträffade	happened	0	0	1	0
legat	formed	0	0	1	0
legat	layed	0	0	1	0
uppbyggnad	construction	0	0	1	1
uppbyggnad	structure	0	0	1	0
storhetstid	heyday	0	0	1	0
liberala	liberal	0	0	1	0
servrar	servers	0	0	1	0
nederländska	netherlands	0	0	1	0
nederländska	dutch	0	0	1	0
domstolar	courts	0	0	1	0
geografi	geography	0	0	1	1
genom	through	0	0	1	1
tyskt	german	0	0	1	0
korrekt	proper	0	0	1	0
korrekt	correct	0	0	1	1
energikällor	energy resources	0	0	1	0
energikällor	energy sources	0	0	1	0
energikällor	sources of energy	0	0	1	0
mandelas	mandelas	0	0	1	0
mandelas	mandela's	0	0	1	0
kollapsade	collapsed	0	0	1	0
närmast	nearest	0	0	1	1
närmast	closest	0	0	1	1
närmast	mediately	0	0	1	0
tyska	german	0	0	1	0
tyske	german	0	0	1	0
tillämpningar	applications	0	0	1	0
tillämpningar	implementations	0	0	1	0
tillämpningar	situations	0	0	1	0
träffar	meets	0	0	1	0
träffar	hits	0	0	1	0
on	on	0	0	1	0
om	of	0	0	1	1
om	for	0	0	1	1
om	if	0	0	1	1
uppdelade	divided	0	0	1	0
indianska	red indian	0	0	1	0
indianska	amerindian	0	0	1	0
indianska	native american	0	0	1	0
träffat	met	0	0	1	0
spelet	the game	0	0	1	0
spelet	game	0	0	1	0
og	og	0	0	1	0
of	of	0	0	1	0
of	av	0	0	1	0
oc	oc	0	0	1	0
oc	o.c.	0	0	1	0
gäst	guest	0	0	1	1
stand	stand	0	0	1	0
framträdanden	the trades of	0	0	1	0
framträdanden	appearances	0	0	1	0
os	os	0	0	1	0
spelen	the games	0	0	1	0
spelen	games	0	0	1	0
koppling	clutch	0	0	1	1
koppling	connection	0	0	1	1
cambridge	cambridge	0	0	1	0
säljs	sold	0	0	1	0
sälja	sell	0	0	1	1
tolkning	interpretations	0	0	1	0
tolkning	interpretation	0	0	1	0
domstol	court	0	0	1	1
burton	burton	0	0	1	0
erövrades	conquered	0	0	1	0
erövrades	(was) conquered	0	0	1	0
erövrades	concoured	0	0	1	0
sfären	spheres	0	0	1	0
sfären	sphere	0	0	1	0
befinna	be	0	0	1	1
upprättade	established	0	0	1	0
upprättade	prepared	0	0	1	0
medlemsstaternas	member	0	0	1	0
medlemsstaternas	member state	0	0	1	0
medlemsstaternas	member states	0	0	1	0
nåddes	reached	0	0	1	0
deltar	participates	0	0	1	0
deltar	part	0	0	1	0
fisk	fish	0	0	1	1
innehöll	contained a ban on	0	0	1	0
innehöll	include	0	0	1	0
innehöll	containing	0	0	1	0
valley	valley	0	0	1	0
serbien	serbia	0	0	1	0
lärt	learned	0	0	1	0
lärt	learnt	0	0	1	0
utgångspunkt	starting point	0	0	1	0
utgångspunkt	point of departure	0	0	1	1
avbröts	canceled	0	0	1	0
avbröts	interrupted	0	0	1	0
flyga	fly	0	0	1	1
inriktning	direction	0	0	1	0
inriktning	orientation	0	0	1	1
inriktning	alignment	0	0	1	1
hävdade	argued	0	0	1	0
hävdade	claimed	0	0	1	0
lära	lara	0	0	1	0
lära	learn	0	0	1	0
lära	get to know	0	0	1	0
ökningen	increase	0	0	1	0
ökningen	the increase	0	0	1	0
ingredienser	ingredients	0	0	1	0
ingredienser	the ingredients	0	0	1	0
ingredienser	ingredient	0	0	1	0
förändra	change; alter; replace	0	0	1	0
förändra	change	0	0	1	1
manuskript	manuscript	0	0	1	1
manuskript	script	0	0	1	1
raúl	raul	0	0	1	0
varning	warning	0	0	1	1
överraskande	surprisingly	0	0	1	0
stövare	beagle	0	0	1	1
stövare	hound	0	0	1	0
chaplin	chaplin	0	0	1	0
kvinnornas	womens	0	0	1	0
kvinnornas	the women's	0	0	1	0
kvinnornas	women	0	0	1	0
taylor	taylor	0	0	1	0
åländska	Åland swedish	0	0	1	0
åländska	aland	0	0	1	0
felix	felix	0	0	1	0
fjorton	fourteen	0	0	1	1
påverkats	influenced	0	0	1	0
påverkats	affected	0	0	1	0
avstå	desist	0	0	1	1
avstå	non	0	0	1	0
avstå	refrain	0	0	1	1
liverpool	liverpool	0	0	1	1
begått	committed	0	0	1	0
begått	comitted	0	0	1	0
bestämd	fixed	0	0	1	1
nämnas	mentioned	0	0	1	0
nämnas	worth mentioning	0	0	1	0
nämnas	include	0	0	1	0
upptäcker	discoveries	0	0	1	0
upptäcker	discover	0	0	1	0
upptäcker	discovers	0	0	1	0
skulder	liabilities	0	0	1	1
skulder	debts	0	0	1	0
skulder	debt	0	0	1	0
kretsen	the order	0	0	1	0
kretsen	circuit	0	0	1	0
roses	roses	0	0	1	0
ovanför	over	0	0	1	1
ovanför	above the	0	0	1	0
ovanför	above	0	0	1	1
utgifter	expenditure	0	0	1	1
utgifter	expenses	0	0	1	0
babylon	babylonia	0	0	1	0
babylon	babylon	0	0	1	0
visade	showed	0	0	1	0
visade	showed; displayed	0	0	1	0
östeuropa	eastern europe	0	0	1	1
östeuropa	east europe	0	0	1	0
separata	separate	0	0	1	0
grupp	group	0	0	1	1
ockupation	occupation	0	0	1	1
gården	farm	0	0	1	0
gården	courtyard; house; farm (-house)	0	0	1	0
gården	garden	0	0	1	0
symbol	symbol	0	0	1	1
missbruk	addiction	0	0	1	1
missbruk	abuse	0	0	1	1
sjätte	sixth	0	0	1	1
vinnaren	winner	0	0	1	0
vinnaren	the winner	0	0	1	0
symtomen	symptoms	0	0	1	0
symtomen	the symptoms	0	0	1	0
symtomen	ymptoms	0	0	1	0
mån	concerned	0	0	1	0
mån	mon	0	0	1	0
villkor	conditions	0	0	1	0
villkor	condition	0	0	1	1
distriktet	district	0	0	1	0
författning	constitution	0	0	1	1
barcelona	barcelona	0	0	1	0
calle	calle	0	0	1	0
erfarenhet	experience	0	0	1	1
visby	visby	0	0	1	0
all	any	0	0	1	1
ali	ali	0	0	1	0
alf	alf	0	0	1	0
separat	seperate	0	0	1	0
separat	separate	0	0	1	1
konsekvens	impact	0	0	1	0
konsekvens	consequence	0	0	1	1
konsekvent	consistent	0	0	1	1
konsekvent	consistency	0	0	1	0
invånare	resident (-s)	0	0	1	0
invånare	inhabitants	0	0	1	0
utomliggande	external; ex-territorial	0	0	1	0
utomliggande	outlying	0	0	1	0
sakrament	sacrament	0	0	1	1
krisen	crisis	0	0	1	0
krisen	the crisis	0	0	1	0
dödsstraff	death penalty	0	0	1	0
förbundet	the union	0	0	1	0
förbundet	association	0	0	1	0
uppdrag	job	0	0	1	0
uppdrag	missions	0	0	1	0
uppdrag	mission	0	0	1	1
persiska	persian	0	0	1	0
funktionerna	functions	0	0	1	0
funktionerna	the functions	0	0	1	0
säsongerna	seasons	0	0	1	0
säsongerna	sason organize	0	0	1	0
kapitulerade	surrendered	0	0	1	0
gary	gary	0	0	1	0
program	application	0	0	1	0
cykeln	there are two meanings in the context - cycle and bicycle	0	0	1	0
cykeln	cycle	0	0	1	0
kvar	left	0	0	1	1
förbundsstat	federal	0	0	1	0
förbundsstat	federal state	0	0	1	1
började	started	0	0	1	0
började	began	0	0	1	0
litet	small	0	0	1	1
solen	the sun	0	0	1	0
solen	sol	0	0	1	0
song	song	0	0	1	0
far	father	0	0	1	1
fas	phase	0	0	1	1
fat	barrel	0	0	1	1
fat	fat	0	0	1	0
runtom	throughout	0	0	1	0
runtom	around	0	0	1	0
simpsons	simpsons	0	0	1	0
högtid	festival	0	0	1	1
högtid	festival; holiday	0	0	1	0
svårigheter	difficulties	0	0	1	0
svårigheter	hardships	0	0	1	0
fan	devil	0	0	1	1
fan	fan	0	0	1	1
sony	sony	0	0	1	0
främja	further	0	0	1	1
främja	promote	0	0	1	1
främja	promoting	0	0	1	0
liten	small	0	0	1	1
unionens	the union	0	0	1	0
unionens	european union	0	0	1	0
unionens	the union's	0	0	1	0
tjeckiska	czech	0	0	1	0
choklad	chocolate	0	0	1	1
knutsson	knutsson	0	0	1	0
nedåt	down	0	0	1	1
nedåt	downward	0	0	1	1
nedåt	down; downwards	0	0	1	0
list	cunning	0	0	1	1
hallucinationer	hallucinations	0	0	1	0
behöll	retained	0	0	1	0
behöll	kept	0	0	1	0
gäng	group	0	0	1	0
gäng	gang	0	0	1	1
gäng	thread	0	0	1	0
konflikt	conflict	0	0	1	1
konflikt	conflict; strife	0	0	1	0
personlighetsstörningar	personality disorders	0	0	1	0
författare	forfatare	0	0	1	0
författare	author	0	0	1	1
lisa	lisa	0	0	1	0
enastående	outstanding	0	0	1	1
enastående	exceptional	0	0	1	0
programme	programme	0	0	1	0
mäktigaste	powerful	0	0	1	0
mäktigaste	most powerful	0	0	1	0
hitta	come up	0	0	1	0
hitta	see	0	0	1	0
hitta	find	0	0	1	1
hitta	make up	0	0	1	0
grekland	greece	0	0	1	1
ted	ted	0	0	1	0
istiden	ice age	0	0	1	0
istiden	the ice age	0	0	1	0
tex	for example	0	0	1	0
tex	e.g.	0	0	1	0
design	design	0	0	1	1
haag	haag	0	0	1	0
haag	the hague	0	0	1	0
kärnvapen	nuclear	0	0	1	0
kärnvapen	nuclear weapons	0	0	1	0
usama	osama	0	0	1	0
usama	usama	0	0	1	0
enklaste	the simplest	0	0	1	0
enklaste	easiest	0	0	1	0
sun	sun	0	0	1	0
vaginalt	vaginal	0	0	1	0
kinesiska	chinese	0	0	1	0
version	version	0	0	1	1
spelning	gig	0	0	1	0
spelning	playing	0	0	1	0
sur	acidic	0	0	1	0
sur	sour	0	0	1	1
guns	guns	0	0	1	0
christian	christian	0	0	1	0
dottern	the daughter	0	0	1	0
dottern	daughter	0	0	1	0
framgången	success	0	0	1	0
framgången	the success	0	0	1	0
regerade	reigned	0	0	1	0
försvaret	the defense	0	0	1	0
försvaret	repository	0	0	1	0
leeds	leeds	0	0	1	0
gång	once	0	0	1	0
gång	time	0	0	1	1
norden	scandinavia; (nordic area; region)	0	0	1	0
norden	the nordic countries	0	0	1	0
norden	north	0	0	1	0
nordens	the scandinavian countries'	0	0	1	0
nordens	scandinavia	0	0	1	0
nordens	nordic	0	0	1	0
folktro	popular belief	0	0	1	0
folktro	folklore	0	0	1	1
soloalbum	solo album	0	0	1	0
säkerhet	safety; security	0	0	1	0
säkerhet	security	0	0	1	1
magnitud	magnitude	0	0	1	1
arabemiraten	united arab emirates	0	0	1	0
arabemiraten	uae	0	0	1	0
arabemiraten	the arab emirate	0	0	1	0
snus	snuff	0	0	1	1
uppkomst	origin	0	0	1	1
uppkomst	onset	0	0	1	0
kategorispelare	category player	0	0	1	0
filmerna	films	0	0	1	0
filmerna	the movies	0	0	1	0
proteinet	protein	0	0	1	0
proteinet	the protein	0	0	1	0
syfte	purpose	0	0	1	0
syfte	view	0	0	1	0
syfta	aim	0	0	1	0
syfta	refer	0	0	1	0
smak	taste	0	0	1	1
smak	flavoring	0	0	1	0
socialdemokraterna	members of the social democracy	0	0	1	0
socialdemokraterna	social democratic	0	0	1	0
anarkism	anarchism	0	0	1	1
anarkism	anarchy	0	0	1	0
ändå	still	0	0	1	1
ändå	spirit	0	0	1	0
branden	fire	0	0	1	0
branden	the fire	0	0	1	0
anc	anc	0	0	1	0
autonom	independent	0	0	1	0
autonom	autonomic	0	0	1	0
besittningar	holdings	0	0	1	0
besittningar	possessions	0	0	1	0
genomsnittliga	average	0	0	1	0
israel	israel	0	0	1	0
israel	israeli	0	0	1	0
permanenta	permanent	0	0	1	0
cellerna	cells	0	0	1	0
cellerna	the cells	0	0	1	0
akademiens	academy	0	0	1	0
akademiens	the academy's	0	0	1	0
akademiens	attend	0	0	1	0
glas	glass	0	0	1	1
anges	mention	0	0	1	0
anges	is put at	0	0	1	0
anges	specified	0	0	1	0
jönköpings	jönköpings	0	0	1	0
jönköpings	jonkopings	0	0	1	0
floyd	floyd	0	0	1	0
livslängd	life	0	0	1	1
livslängd	life expectancy	0	0	1	0
glad	happy	0	0	1	1
naturligt	natural	0	0	1	0
legender	legends	0	0	1	0
salvador	salvador	0	0	1	0
decenniet	decade	0	0	1	0
decennier	decades	0	0	1	0
kryddor	spices	0	0	1	0
mussolini	mussolini	0	0	1	0
mussolini	mossolini	0	0	1	0
kommendör	commandor	0	0	1	0
kommendör	commander	0	0	1	1
pony	pony	0	0	1	0
brown	brown	0	0	1	0
grundläggande	because lag of	0	0	1	0
grundläggande	primary	0	0	1	0
grundläggande	fundamental	0	0	1	1
duett	duet	0	0	1	1
bosatt	resident	0	0	1	1
bosatt	lived	0	0	1	0
årets	the year's	0	0	1	0
årets	this year's	0	0	1	0
årets	year	0	0	1	0
huvudort	main town	0	0	1	0
huvudort	principal town	0	0	1	0
jordens	earth	0	0	1	0
elektrisk	electric	0	0	1	1
elektrisk	elektirsk	0	0	1	0
historiskt	historic	0	0	1	0
historiskt	historically	0	0	1	0
historiskt	historical	0	0	1	0
court	court	0	0	1	0
breaking	breakingpoint	0	0	1	0
breaking	breaking	0	0	1	0
genomsnittet	average	0	0	1	0
genomsnittet	the average	0	0	1	0
brittisk	british	0	0	1	1
satanism	satanism	0	0	1	0
satanism	satanic	0	0	1	0
historiska	historical	0	0	1	0
ihåg	remember	0	0	1	0
skolan	school	0	0	1	0
indelade	divided	0	0	1	0
indelade	divided into	0	0	1	0
fört	led	0	0	1	0
fört	lead	0	0	1	0
förr	sooner; past	0	0	1	0
förr	sooner	0	0	1	1
förr	before	0	0	1	1
förs	rapids	0	0	1	0
förs	led	0	0	1	0
förs	out	0	0	1	0
taget	a time (practically; virtually; any; at all)	0	0	1	0
taget	time	0	0	1	0
årligen	annually	0	0	1	1
årligen	yearly	0	0	1	1
årligen	annual	0	0	1	0
sven	sven	0	0	1	0
tagen	taken	0	0	1	1
producerad	produced	0	0	1	0
före	before	0	0	1	1
före	present	0	0	1	0
före	ahead (of)	0	0	1	0
föra	pre	0	0	1	0
föra	lead	0	0	1	1
atomer	atoms	0	0	1	0
regnar	rains	0	0	1	0
regnar	raining	0	0	1	0
fördelen	advantage	0	0	1	0
fördelen	the advantage	0	0	1	0
anarkistiska	anarchistic	0	0	1	0
anarkistiska	anarchist	0	0	1	0
praktiska	practical	0	0	1	0
frågorna	questions	0	0	1	0
frågorna	questions; issues	0	0	1	0
bildade	formed	0	0	1	0
vänster	left	0	0	1	1
därav	thereof	0	0	1	0
praktiskt	convenient	0	0	1	0
homosexuella	homosexual	0	0	1	0
homosexuella	gay	0	0	1	0
grande	grande	0	0	1	0
grande	grand	0	0	1	0
moraliska	moral	0	0	1	0
greklands	greek gloss	0	0	1	0
greklands	greek country	0	0	1	0
greklands	greece's	0	0	1	0
friidrott	athletics	0	0	1	1
friidrott	track and field	0	0	1	0
avvisade	rejected	0	0	1	0
september	september	0	0	1	1
emmanuel	emmanuel	0	0	1	0
mission	mission	0	0	1	1
australien	australian	0	0	1	0
australien	australia	0	0	1	1
retoriska	rhetorical	0	0	1	0
självständiga	independent	0	0	1	0
självständiga	sjalvstandiga	0	0	1	0
närstående	relative	0	0	1	0
närstående	relatives	0	0	1	0
närstående	kindred	0	0	1	0
islam	islam	0	0	1	1
lyder	reads	0	0	1	0
lyder	obeys	0	0	1	0
rika	rich	0	0	1	0
abbey	abbey	0	0	1	0
ärftliga	genetic	0	0	1	0
rikt	target	0	0	1	0
rikt	rich	0	0	1	0
prag	prague	0	0	1	1
stephen	stephen	0	0	1	0
argentina	argentina	0	0	1	1
fenomenet	the phenomenon	0	0	1	0
fenomenet	phenomenon	0	0	1	0
kategorieuropeiska	european category	0	0	1	0
kategorieuropeiska	europe category	0	0	1	0
styret	gate	0	0	1	0
medborgerliga	civil	0	0	1	0
genomgående	consistently	0	0	1	0
genomgående	through	0	0	1	1
genomgående	pervading	0	0	1	1
postumt	posthumous award	0	0	1	0
postumt	posthumously	0	0	1	0
chicago	chicago	0	0	1	1
landborgen	the ridge	0	0	1	0
marcus	marcus	0	0	1	0
skönlitteratur	nonfiction	0	0	1	0
skönlitteratur	fiction	0	0	1	1
journalisten	journalist	0	0	1	0
journalisten	the journalist	0	0	1	0
forna	former	0	0	1	0
forna	previous	0	0	1	0
stilen	style	0	0	1	0
viktigt	important	0	0	1	0
slidan	the vagina	0	0	1	0
slidan	vagina	0	0	1	0
slidan	vaginal	0	0	1	0
journalister	journalists	0	0	1	0
principer	principals	0	0	1	0
principer	principles	0	0	1	0
kustlinje	coastline	0	0	1	1
ringar	rings	0	0	1	0
drycken	beverage	0	0	1	0
drycken	the drink	0	0	1	0
betyg	grades	0	0	1	0
betyg	marks	0	0	1	0
brother	brother	0	0	1	0
århundraden	centuries	0	0	1	0
aldrig	never	0	0	1	1
mongoliet	mongolia	0	0	1	0
stenar	stones	0	0	1	0
stenar	blocks	0	0	1	0
beyoncé	beyoncé	0	0	1	0
beyoncé	beyoncè	0	0	1	0
beyoncé	beyonce	0	0	1	0
ollonet	penis head	0	0	1	0
ollonet	glans	0	0	1	0
ollonet	the glans	0	0	1	0
förhistorisk	forhistorisk	0	0	1	0
förhistorisk	prehistorian	0	0	1	0
nepal	nepal	0	0	1	1
europas	europe	0	0	1	0
hill	hill	0	0	1	0
delstat	state	0	0	1	0
delstat	land	0	0	1	0
arvid	arvid	0	0	1	0
benjamin	benjamin	0	0	1	0
poliser	police (-men; -women)	0	0	1	0
poliser	police	0	0	1	0
återvände	returned	0	0	1	0
återvände	returning	0	0	1	0
väldigt	very	0	0	1	1
islamistiska	islamic	0	0	1	0
islamistiska	islamist	0	0	1	0
densiteten	density	0	0	1	0
rörande	on	0	0	1	0
rörande	concerning	0	0	1	1
statsöverhuvud	head of state	0	0	1	0
översatt	translated	0	0	1	0
översatt	the translation	0	0	1	0
avsett	avset	0	0	1	0
avsett	regard	0	0	1	0
avsett	intended	0	0	1	0
förtroende	confidence	0	0	1	1
förtroende	trust	0	0	1	1
kritiserat	criticized	0	0	1	0
kritiserat	criticised	0	0	1	0
väldiga	immense	0	0	1	0
väldiga	mighty	0	0	1	0
väldiga	vast	0	0	1	0
spelades	filmed	0	0	1	0
kritiserar	criticize	0	0	1	0
polisen	police	0	0	1	0
polisen	the police	0	0	1	0
faller	fall	0	0	1	0
fallet	case	0	0	1	0
fallet	the case	0	0	1	0
stavningen	spelling	0	0	1	0
stavningen	the spelling	0	0	1	0
konsumtionen	the consumtion	0	0	1	0
konsumtionen	consumption	0	0	1	0
bekräftade	confirmed	0	0	1	0
pendeltåg	commuter train	0	0	1	0
pendeltåg	commuter	0	0	1	0
soundtrack	soundtrack	0	0	1	0
soundtrack	sound rack	0	0	1	0
fallen	case	0	0	1	0
fallen	cases	0	0	1	0
sträckan	distance	0	0	1	0
sträckan	the distance	0	0	1	0
sår	sir	0	0	1	0
sår	wound	0	0	1	1
aminosyror	aminosynor	0	0	1	0
aminosyror	amino acids	0	0	1	0
såg	see	0	0	1	0
såg	saw	0	0	1	1
filosofins	philosophy	0	0	1	0
filosofins	the philosophy	0	0	1	0
colombia	colombia	0	0	1	1
pablo	pablo	0	0	1	0
bland	blamd	0	0	1	0
bland	inter	0	0	1	0
bland	including	0	0	1	0
äldsta	oldest	0	0	1	0
blanc	blanc	0	0	1	0
story	story	0	0	1	1
spred	spread	0	0	1	0
automobile	automobile	0	0	1	0
misslyckas	fail	0	0	1	1
misslyckas	fails	0	0	1	0
stort	large	0	0	1	0
stort	big	0	0	1	0
motiveringen	the motivation	0	0	1	0
motiveringen	ground	0	0	1	0
storm	storm	0	0	1	1
kristendomens	christianity	0	0	1	0
kristendomens	the christianity's	0	0	1	0
kristendomens	christianity's	0	0	1	0
stora	large	0	0	1	0
stora	big	0	0	1	0
ecuador	ecuador	0	0	1	1
familjerna	families	0	0	1	0
mikael	mikael	0	0	1	0
minoritetsspråk	minority language	0	0	1	0
minoritetsspråk	minority	0	0	1	0
hotel	hotel	0	0	1	0
böcker	useful downloads archive	0	0	1	0
böcker	books	0	0	1	1
kongress	congress	0	0	1	1
serotonin	serotonin	0	0	1	0
framtiden	future	0	0	1	0
framtiden	the future	0	0	1	0
hotet	threat	0	0	1	0
hotet	the threat	0	0	1	0
hotet	the threath	0	0	1	0
fattigaste	the poorest	0	0	1	0
fattigaste	poorest	0	0	1	0
siffra	number	0	0	1	0
siffra	figure	0	0	1	1
king	king	0	0	1	0
illegala	illegal	0	0	1	0
illegala	irregular	0	0	1	0
matcherna	the games	0	0	1	0
matcherna	games	0	0	1	0
smält	melted	0	0	1	0
kina	china	0	0	1	1
röda	red	0	0	1	0
dans	dance	0	0	1	1
guden	god	0	0	1	0
guden	the god	0	0	1	0
kategorin	category	0	0	1	0
kategorin	the category	0	0	1	0
klubb	club	0	0	1	1
filosofin	philosophy	0	0	1	0
filosofin	the philosophy	0	0	1	0
kusin	cousin	0	0	1	1
tilldelas	assigned	0	0	1	0
tilldelas	award	0	0	1	0
föreligger	is	0	0	1	0
föreligger	exist	0	0	1	0
tabell	table	0	0	1	1
tabell	chart	0	0	1	1
tabell	tabel	0	0	1	0
humör	temper	0	0	1	1
humör	mood	0	0	1	1
divisionen	division	0	0	1	0
wilson	wilson	0	0	1	0
bedriver	manage	0	0	1	0
bedriver	conducts	0	0	1	0
bedriver	operate	0	0	1	0
inriktningar	direction	0	0	1	0
inriktningar	specializations	0	0	1	0
dialekt	dialect	0	0	1	1
dialekt	brogue	0	0	1	0
överenskommelse	deal	0	0	1	1
överenskommelse	arrangement	0	0	1	0
judas	judas	0	0	1	1
unge	young	0	0	1	1
unge	kid	0	0	1	1
folkgrupper	communities	0	0	1	0
folkgrupper	ethnic groups	0	0	1	0
electric	electic	0	0	1	0
electric	electric	0	0	1	0
dagliga	daily	0	0	1	0
park	park	0	0	1	1
lätt	easy	0	0	1	1
naturvetenskapliga	science	0	0	1	0
naturvetenskapliga	scientific	0	0	1	0
dagligt	daily	0	0	1	0
industrialiserade	industrialized	0	0	1	0
skräck	fear	0	0	1	0
skräck	horror	0	0	1	1
mineral	minerals	0	0	1	0
mineral	mineral	0	0	1	1
windows	windows	0	0	1	0
medelhavsområdet	the mediterranean region	0	0	1	0
medelhavsområdet	mediterranean	0	0	1	0
medelhavsområdet	the mediterranean area	0	0	1	0
influensan	the influenza	0	0	1	0
influensan	flu	0	0	1	0
statsskick	polity	0	0	1	0
statsskick	form of government	0	0	1	0
statsskick	government	0	0	1	1
osäkert	insecure	0	0	1	0
osäkert	unclear	0	0	1	0
osäkert	uncertain	0	0	1	0
kosovo	kosovo	0	0	1	0
tjugo	twenty	0	0	1	1
växjö	vaxjo	0	0	1	0
växjö	växjö	0	0	1	0
ursprungliga	original	0	0	1	0
kolonialism	colonialism	0	0	1	1
allmän	allman	0	0	1	0
allmän	general	0	0	1	1
tilly	tilly	0	0	1	0
tills	until the	0	0	1	0
tills	until	0	0	1	1
agnosticism	agnosticism	0	0	1	1
canaria	canaria	0	0	1	0
grace	grace	0	0	1	1
känsliga	susceptible	0	0	1	0
känsliga	1st&2nd: fragile 3rd: sensitive	0	0	1	0
känsliga	bilge accordance	0	0	1	0
moses	moses	0	0	1	0
his	his	0	0	1	0
hit	to here	0	0	1	0
hit	here	0	0	1	1
försöken	trials	0	0	1	0
försöken	attempts	0	0	1	0
försöken	the tries	0	0	1	0
hiv	hiv	0	0	1	0
märta	märta	0	0	1	0
stormakterna	great powers	0	0	1	0
inklusive	including	0	0	1	1
vardera	either	0	0	1	1
vardera	each	0	0	1	1
b	b	0	0	1	0
jobbade	worked	0	0	1	0
försöker	try	0	0	1	0
försöker	tries	0	0	1	0
försöker	trying	0	0	1	0
sofie	sofie	0	0	1	0
solsystemet	the solar system	0	0	1	0
solsystemet	solar system`	0	0	1	0
budapest	budapest	0	0	1	0
utvidgade	expanded	0	0	1	0
tvkanaler	tv-channels	0	0	1	0
tvkanaler	tv channels	0	0	1	0
mediciner	medicines	0	0	1	0
avtal	agreement; deal	0	0	1	0
avtal	agreement	0	0	1	1
avtal	contract	0	0	1	1
tidszon	timezone	0	0	1	0
tidszon	time zone	0	0	1	0
vincent	vincent	0	0	1	0
virginia	virginia	0	0	1	1
reagan	reagan	0	0	1	0
utsatt	exposed	0	0	1	1
bars	bar	0	0	1	0
bars	carried	0	0	1	0
etiopien	ethiopia	0	0	1	1
etiopien	ethiopian	0	0	1	0
art	kind	0	0	1	1
art	art	0	0	1	0
bart	offense	0	0	1	0
bart	bart	0	0	1	0
arv	heritage	0	0	1	1
fiske	fishing	0	0	1	1
dödsorsaken	cause of death	0	0	1	0
möta	meet	0	0	1	1
möta	face	0	0	1	0
möte	meeting	0	0	1	1
are	are	0	0	1	0
arg	angry	0	0	1	1
flyttade	moved	0	0	1	0
arm	arm	0	0	1	1
barn	child	0	0	1	1
bortsett	except	0	0	1	0
bortsett	apart	0	0	1	0
planeras	is planned	0	0	1	0
planeras	planned	0	0	1	0
planerar	is planning	0	0	1	0
planerar	plan	0	0	1	0
planerar	planned	0	0	1	0
uppskatta	estimate	0	0	1	1
uppskatta	appreciate	0	0	1	1
inga	not	0	0	1	0
inga	no	0	0	1	1
rod	rod	0	0	1	0
planerat	planned	0	0	1	0
invaldes	elected	0	0	1	0
invaldes	was elected	0	0	1	0
hårdvara	hardware	0	0	1	1
hårdvara	hardwere	0	0	1	0
källor	source	0	0	1	0
källor	calla lilies	0	0	1	0
växthuseffekten	the greenhouse effect	0	0	1	0
växthuseffekten	greenhouse effect	0	0	1	0
nätverk	network	0	0	1	1
law	law	0	0	1	0
planerad	planned	0	0	1	0
muslim	muslim	0	0	1	1
fördelas	be allocated	0	0	1	0
fördelas	distribute	0	0	1	0
fördelas	distributed	0	0	1	0
ändras	be changed	0	0	1	0
ändras	change	0	0	1	0
såväl	both	0	0	1	0
såväl	as well as	0	0	1	0
vände	reversed	0	0	1	0
vände	turned	0	0	1	0
vända	turn	0	0	1	1
vända	habituated	0	0	1	0
herrar	gentlemen	0	0	1	0
herrar	men	0	0	1	0
uppkom	arose	0	0	1	0
kämpade	decreased	0	0	1	0
kämpade	fought	0	0	1	0
uppträder	appears	0	0	1	0
uppträder	performs	0	0	1	0
uppträder	occur	0	0	1	0
tiderna	the times	0	0	1	0
tiderna	time	0	0	1	0
tiderna	ages	0	0	1	0
tiderna	times	0	0	1	0
startades	started	0	0	1	0
operan	opera	0	0	1	0
operan	the opera	0	0	1	0
roman	novel	0	0	1	1
öarna	the islands	0	0	1	0
öarna	islands	0	0	1	0
hypotesen	the hypothesis	0	0	1	0
hypotesen	hypothesis	0	0	1	0
görs	is	0	0	1	0
görs	made	0	0	1	0
görs	is made to	0	0	1	0
borta	gone	0	0	1	1
borta	away	0	0	1	1
räknar	counts	0	0	1	0
räknar	counter	0	0	1	0
vidare	moreover	0	0	1	0
vidare	furthermore	0	0	1	1
vidare	further	0	0	1	1
räknat	calculated	0	0	1	0
räknat	counted	0	0	1	0
göra	do	0	0	1	1
göra	do; doing	0	0	1	0
nationalpark	national park	0	0	1	0
besegrade	defeated	0	0	1	0
tränare	coach	0	0	1	1
tränare	tranae	0	0	1	0
hypoteser	hypotheses	0	0	1	0
hypoteser	hypothesis	0	0	1	0
gäster	guests	0	0	1	0
ps	ps	0	0	1	0
ps	p.s	0	0	1	0
ps	p.s.	0	0	1	0
java	java	0	0	1	1
skrev	said	0	0	1	0
personalen	personnel	0	0	1	0
personalen	the staff	0	0	1	0
nationalförsamlingen	nationaforsamlingen	0	0	1	0
nationalförsamlingen	national assembly	0	0	1	0
kungafamiljen	the royal family	0	0	1	0
johannes	johannes	0	0	1	0
johannes	john	0	0	1	0
pc	pc	0	0	1	0
pc	personal computer	0	0	1	0
karriären	career	0	0	1	0
karriären	the career	0	0	1	0
byxor	pants	0	0	1	1
ska	will	0	0	1	0
ska	shall	0	0	1	0
ph	ph	0	0	1	0
pi	pi	0	0	1	1
chandler	chandler	0	0	1	0
flight	flights	0	0	1	0
flight	flight	0	0	1	0
småningom	when the time comes	0	0	1	0
småningom	eventually	0	0	1	0
togs	taken	0	0	1	0
togs	were taken	0	0	1	0
publiken	the audience	0	0	1	0
publiken	audience	0	0	1	0
sydafrikas	of south africa	0	0	1	0
sydafrikas	south african	0	0	1	0
sydafrikas	south africa's	0	0	1	0
passade	suiting	0	0	1	0
passade	suited	0	0	1	0
passade	fit; suited	0	0	1	0
konflikter	conflicts	0	0	1	0
konflikter	conflict	0	0	1	0
konflikten	the conflict	0	0	1	0
konflikten	conflict	0	0	1	0
deltog	participated	0	0	1	0
medelålder	middle age	0	0	1	1
medelålder	mean age	0	0	1	0
inspelningar	recordings	0	0	1	0
styr	controls	0	0	1	0
ris	rice	0	0	1	1
effektiv	effective	0	0	1	1
rik	rich	0	0	1	1
rik	rish	0	0	1	0
fullständig	full	0	0	1	1
fullständig	complete	0	0	1	1
fullständig	n/a	0	0	1	0
spåra	track	0	0	1	1
spåra	trace	0	0	1	1
byggnaderna	building	0	0	1	0
byggnaderna	buildings	0	0	1	0
byggnaderna	the buildings	0	0	1	0
skeppen	the ships	0	0	1	0
fysisk	natural	0	0	1	0
fysisk	physical	0	0	1	1
demografi	demographics	0	0	1	0
demografi	demography	0	0	1	1
tidpunkten	the time	0	0	1	0
tidpunkten	the moment	0	0	1	0
tidpunkten	time	0	0	1	0
ideologier	ideologies	0	0	1	0
sjunkit	decreased	0	0	1	0
bortgång	passing	0	0	1	1
bortgång	death	0	0	1	1
på	on	0	0	1	1
på	at	0	0	1	1
på	in	0	0	1	1
omgivning	surrounding	0	0	1	0
omgivning	surroundings	0	0	1	0
omgivning	ambient	0	0	1	0
järnvägarna	the railways	0	0	1	0
järnvägarna	railways	0	0	1	0
spears	spears	0	0	1	0
skeppet	the ship	0	0	1	0
skeppet	nave	0	0	1	0
byar	villages	0	0	1	0
uppbyggd	structured	0	0	1	0
uppbyggd	structered	0	0	1	0
uppbyggd	built-up	0	0	1	0
förklarar	explain	0	0	1	0
förklarar	explains	0	0	1	0
uppbyggt	structured	0	0	1	0
gräs	grass	0	0	1	1
kokpunkt	having a boiling point	0	0	1	0
kokpunkt	boiling point	0	0	1	0
vinklar	angle	0	0	1	0
vinklar	angles	0	0	1	0
finansiera	fund	0	0	1	0
finansiera	finance	0	0	1	1
italiensk	italian	0	0	1	1
sjunga	access	0	0	1	0
sjunga	sing	0	0	1	1
edge	edge	0	0	1	0
utnämndes	was declared	0	0	1	0
utnämndes	appointed	0	0	1	0
vetenskapen	the science	0	0	1	0
vetenskapen	science	0	0	1	0
kyrkans	the churche's	0	0	1	0
kyrkans	the church's	0	0	1	0
kyrkans	church	0	0	1	0
alfabet	alphabets	0	0	1	0
alfabet	alphabet	0	0	1	1
fängslade	inprisoned	0	0	1	0
fängslade	confine	0	0	1	0
fängslade	imprisoned	0	0	1	0
bokstäver	letters	0	0	1	0
kontinentala	continental	0	0	1	0
reagera	reacting	0	0	1	0
reagera	reaching	0	0	1	0
komplett	complete	0	0	1	1
konstitution	constitution	0	0	1	1
infrastruktur	infrastructure	0	0	1	1
änglar	angels	0	0	1	0
förening	union	0	0	1	1
förening	compound	0	0	1	1
remmer	remmer	0	0	1	0
prince	prince	0	0	1	0
namnet	name	0	0	1	0
namnet	the name	0	0	1	0
winnerbäck	winnerback	0	0	1	0
winnerbäck	winnerbäck	0	0	1	0
skalv	shock	0	0	1	0
skalv	quake	0	0	1	1
minoriteter	minorities	0	0	1	0
bostad	lodge	0	0	1	0
bostad	property	0	0	1	0
omedelbar	instant	0	0	1	1
omedelbar	immediate	0	0	1	1
skall	is	0	0	1	0
skall	shall	0	0	1	1
centralasien	central asia	0	0	1	0
namnen	the names	0	0	1	0
namnen	names	0	0	1	0
namnen	name	0	0	1	0
px|centrerad	px | centric	0	0	1	0
rörelsens	movement	0	0	1	0
rörelsens	operating	0	0	1	0
rörelsens	movements	0	0	1	0
skala	scale	0	0	1	1
skala	scale; size	0	0	1	0
undersöka	study	0	0	1	0
undersöka	understand	0	0	1	0
undersöka	research	0	0	1	0
synnerhet	specially	0	0	1	0
synnerhet	particular	0	0	1	0
djupare	depth	0	0	1	0
djupare	deeper	0	0	1	0
ökad	increase	0	0	1	0
ökad	increased	0	0	1	0
österrike	austria	0	0	1	1
bioetik		1	0	1	0
bioetik	warrior	1	0	1	0
bioetik	bioethics	1	1	0	0
bioetik	wars	1	0	1	0
bioetik	biotik	1	0	1	0
bioetik	bioethic	1	1	0	0
bioetik	bio ethics	1	0	1	0
rastafarianerna	the rastafarian	0	0	1	0
rastafarianerna	rest are faria	0	0	1	0
rastafarianerna	n/a	0	0	1	0
ökar	increasing frequency of	0	0	1	0
ökar	increases	0	0	1	0
begravdes	buried	0	0	1	0
stoppade	stop	0	0	1	0
stoppade	stopped	0	0	1	0
upplevelse	experience	0	0	1	1
exakt	precise	0	0	1	1
exakt	accurately	0	0	1	0
dåvarande	then	0	0	1	1
dåvarande	formerly	0	0	1	0
djävulen	devil	0	0	1	0
djävulen	the devil	0	0	1	0
öster	east	0	0	1	1
guvernör	governor	0	0	1	1
banbrytande	groundbreaking	0	0	1	1
hittar	found	0	0	1	0
hittar	finds	0	0	1	0
hittas	found	0	0	1	0
hittas	be found	0	0	1	0
hittat	found	0	0	1	0
minskning	decline	0	0	1	1
minskning	reduction	0	0	1	1
minskning	decrease	0	0	1	1
landskommun	rural municipality	0	0	1	0
havsnivån	sea level	0	0	1	0
norrut	north	0	0	1	0
bör	live	0	0	1	0
bör	should	0	0	1	0
kongo	congo	0	0	1	1
kongo	kongo	0	0	1	0
lettland	latvia	0	0	1	1
trummis	drummer	0	0	1	0
trummis	trummis	0	0	1	0
begränsade	restricted	0	0	1	0
begränsade	limiting	0	0	1	0
global	global	0	0	1	1
flottan	the fleet	0	0	1	0
flottan	navy	0	0	1	0
flottan	the navy	0	0	1	0
interna	internal	0	0	1	0
håll	ways	0	0	1	0
håll	hold	0	0	1	1
bön	nests	0	0	1	0
bön	prayer	0	0	1	1
grekerna	greeks	0	0	1	0
grekerna	greek	0	0	1	0
ersättning	pay	0	0	1	0
ersättning	remuneration	0	0	1	1
ersättning	replacement	0	0	1	1
prov	test	0	0	1	1
prov	tests	0	0	1	0
fungera	act	0	0	1	0
anne	anne	0	0	1	0
trinidad	trinidad	0	0	1	0
anna	anna	0	0	1	0
turism	tourism	0	0	1	1
diamant	diamond	0	0	1	1
palmes	palme	0	0	1	0
palmes	palme's	0	0	1	0
palmes	plame's	0	0	1	0
producent	prodcuer	1	1	0	0
producent	producer	1	1	1	1
producent	producent; tillverkare	1	0	1	0
producent	producers	1	0	1	0
producent	produce	1	0	1	0
producent	pregnancy	1	0	1	0
anklagades	accused	0	0	1	0
återgick	returned	0	0	1	0
återgick	returning	0	0	1	0
bayern	bavaria	0	0	1	0
bayern	bayern	0	0	1	0
judendom	judaism	0	0	1	1
judendom	jewism	0	0	1	0
kostnaderna	costs	0	0	1	0
kostnaderna	the costs	0	0	1	0
russell	russell	0	0	1	0
russell	rusell	0	0	1	0
virus	virus	0	0	1	1
page	page	0	0	1	1
ande	of	0	0	1	0
ande	spirit	0	0	1	1
dialog	dialogue	0	0	1	1
fotboll	football	0	0	1	1
socialistisk	socialistic	0	0	1	1
socialistisk	socialist	0	0	1	1
oktoberrevolutionen	the october revolution	0	0	1	0
oktoberrevolutionen	october revolution	0	0	1	0
dahléns	dahlens	0	0	1	0
dahléns	dahlen	0	0	1	0
dahléns	dahlén's	0	0	1	0
medborgarna	the citizens	0	0	1	0
medborgarna	citizens	0	0	1	0
reglerna	rules	0	0	1	0
reglerna	rules; regulations	0	0	1	0
svenskspråkiga	swedish speaking	0	0	1	0
svenskspråkiga	swedish-speaking	0	0	1	0
abbas	abbas	0	0	1	0
laget	the team	0	0	1	0
laget	stroke	0	0	1	0
året	the year	0	0	1	0
året	all year	0	0	1	0
året	years	0	0	1	0
dricka	drinking	0	0	1	0
dricka	drink	0	0	1	1
mängder	amounts	0	0	1	0
mängder	amount	0	0	1	0
long	long	0	0	1	0
long	longitude	0	0	1	0
jugoslavien	yugoslavia	0	0	1	1
bagge	bagge	0	0	1	0
bagge	ram	0	0	1	1
bruk	using	0	0	1	0
bruk	use	0	0	1	1
laila	laila	0	0	1	0
sångerska	songstress	0	0	1	0
sångerska	singer	0	0	1	1
ateister	atheists	0	0	1	0
ateister	steister	0	0	1	0
åren	the years	0	0	1	0
åren	years	0	0	1	0
värdefulla	valueable	0	0	1	0
värdefulla	value	0	0	1	0
värdefulla	valuable	0	0	1	0
avslutade	ended	0	0	1	0
avslutade	finished	0	0	1	0
delning	division	0	0	1	1
delning	pitch	0	0	1	0
rasade	collapsed	0	0	1	0
regionen	the region	0	0	1	0
regionen	region	0	0	1	0
dalí	dali	0	0	1	0
kubas	cuba's	0	0	1	0
kubas	cuba	0	0	1	0
hjärta	heart	0	0	1	1
kritikerna	critics	0	0	1	0
kritikerna	the critics	0	0	1	0
kritikerna	critiques	0	0	1	0
delta	delta	0	0	1	1
delta	participate	0	0	1	1
regioner	regions	0	0	1	0
junior	junior	0	0	1	1
medeltidens	ages	0	0	1	0
medeltidens	medieval	0	0	1	0
å	on	0	0	1	0
å	river	0	0	1	1
å	of the	0	0	1	0
planeternas	the planets'	0	0	1	0
planeternas	planets	0	0	1	0
planeternas	the planets	0	0	1	0
styrande	rulers	0	0	1	0
styrande	governing	0	0	1	1
köln	cologne	0	0	1	1
köln	köln	0	0	1	0
homo	homo	0	0	1	0
homo	gay	0	0	1	0
avsevärt	substantially	0	0	1	0
avsevärt	considerably	0	0	1	0
guyana	guyana (name)	0	0	1	0
guyana	guyana	0	0	1	0
tolka	interpreting	0	0	1	0
tolka	interpret	0	0	1	1
fick	got	0	0	1	0
fick	was	0	0	1	0
försvarade	rapid lasted	0	0	1	0
försvarade	defended	0	0	1	0
z	z	0	0	1	0
distinkt	distinct	0	0	1	1
distinkt	distinctive	0	0	1	0
tidens	time's	0	0	1	0
tidens	time	0	0	1	0
tidens	that time's	0	0	1	0
län	state	0	0	1	0
län	between	0	0	1	0
singlarna	singles	0	0	1	0
singlarna	the singles	0	0	1	0
singlarna	simglama	0	0	1	0
tidpunkt	date	0	0	1	1
tidpunkt	time	0	0	1	1
sträckor	distances	0	0	1	0
home	home	0	0	1	0
intressanta	interesting	0	0	1	0
intressanta	of interest	0	0	1	0
graham	graham	0	0	1	0
därutöver	in addition	0	0	1	0
därutöver	addition	0	0	1	0
därutöver	moreover	0	0	1	0
veckorna	weeks	0	0	1	0
rainbow	rainbow	0	0	1	0
stadion	stadium	0	0	1	1
stadion	the stadium	0	0	1	0
vattenånga	steam	0	0	1	1
vattenånga	water vapour	0	0	1	0
psykoterapi	psychotherapy	0	0	1	0
psykoterapi	treatment	0	0	1	0
hanen	the cock	0	0	1	0
hanen	the male	0	0	1	0
hanen	male	0	0	1	0
uppmärksamhet	attention	0	0	1	1
uppmärksamhet	attantion	0	0	1	0
urval	selection	0	0	1	1
skyddas	skyas	0	0	1	0
skyddas	protected	0	0	1	0
skyddas	(is/are) protected	0	0	1	0
skyddar	protection	0	0	1	0
skyddar	protects	0	0	1	0
sutra	sutra	0	0	1	0
feodala	feudal	0	0	1	0
tittarna	the viewers	0	0	1	0
tittarna	viewers	0	0	1	0
medina	medina	0	0	1	0
konvertera	conversion	0	0	1	0
konvertera	convert	0	0	1	1
betyder	means	0	0	1	0
organisk	organic	0	0	1	1
kaspiska	caspian	0	0	1	0
modernismen	modernism	0	0	1	0
klubbens	club	0	0	1	0
vice	vice	0	0	1	0
släppt	self-indulgent	0	0	1	0
släppt	released	0	0	1	0
släppt	relinquished	0	0	1	0
europeiska	european	0	0	1	0
microsoft	microsoft	0	0	1	0
nasa	nasa	0	0	1	0
karma	karma	0	0	1	1
lagstiftning	law-making	0	0	1	0
lagstiftning	regulation	0	0	1	0
europeiskt	europeiskt	0	0	1	0
europeiskt	european	0	0	1	0
nash	' nash	0	0	1	0
nash	nash	0	0	1	0
släppa	release	0	0	1	1
släppa	relaxed	0	0	1	0
psykologi	psychology	0	0	1	1
atombomberna	atom bombs	0	0	1	0
atombomberna	the nuclear bombs	0	0	1	0
atombomberna	atomic bomb	0	0	1	0
tänkandet	thinking	0	0	1	0
tänkandet	the way of thinking	0	0	1	0
tävla	compete	0	0	1	1
kanal	channel	0	0	1	1
mördade	murdered	0	0	1	0
steve	steve	0	0	1	0
jimi	jimi	0	0	1	0
underlättar	make it easier	0	0	1	0
underlättar	facilitates	0	0	1	0
moseboken	genesis	0	0	1	0
kolonialismen	the colonialism	0	0	1	0
kolonialismen	colonialism	0	0	1	0
simon	simon	0	0	1	0
uppmaning	call	0	0	1	0
uppmaning	call; injunction	0	0	1	0
uppmaning	exhortation	0	0	1	1
fortfarande	still	0	0	1	1
romerna	roma	0	0	1	0
romerna	the romani	0	0	1	0
romerna	the romani people	0	0	1	0
uppnå	achieving	0	0	1	0
uppnå	achieve	0	0	1	1
stärkte	strengthened	0	0	1	0
stärkte	increased	0	0	1	0
generellt	generally	0	0	1	1
översvämningar	flooding	0	0	1	0
översvämningar	floodings	0	0	1	0
generella	overall	0	0	1	0
generella	general	0	0	1	0
hinduism	hinduism	0	0	1	1
fotnoter	footnotes	0	0	1	0
pengarna	the money	0	0	1	0
pengarna	money	0	0	1	0
varierar	varies	0	0	1	0
varierar	vary	0	0	1	0
vapen	weapons	0	0	1	0
vapen	weapon	0	0	1	1
kategoritvseriestarter	category television series starts	0	0	1	0
georgien	georgia	0	0	1	1
mesopotamien	mesopotamia	0	0	1	0
sjukdomar	diseases	0	0	1	0
sjukdomar	disease	0	0	1	0
ständig	constant	0	0	1	0
avslutas	close	0	0	1	1
avslutas	ends	0	0	1	0
avslutas	closing	0	0	1	0
avslutat	completed	0	0	1	0
avslutat	finished	0	0	1	0
tvinga	force	0	0	1	1
säkra	reliable	0	0	1	0
säkra	safe	0	0	1	0
säkra	secure	0	0	1	1
historikern	historian	0	0	1	0
historikern	the historian	0	0	1	0
georgier	about	1	0	1	0
georgier	georgian	1	1	0	1
georgier	approximate	1	0	1	0
georgier	the georgians	1	0	1	0
georgier	georgier	1	0	1	0
georgier	georgians	1	1	0	0
lämningar	remains	0	0	1	0
lämningar	remnants	0	0	1	1
anslöt	joined	0	0	1	0
begränsningar	limitations	0	0	1	0
begränsningar	limits	0	0	1	0
demokratiskt	democratic	0	0	1	0
byggt	building	0	0	1	0
byggt	built	0	0	1	0
noter	notes	0	0	1	0
noter	notation	0	0	1	0
ifrågasatt	question	0	0	1	0
ifrågasatt	questioned	0	0	1	0
byggs	building	0	0	1	0
byggs	under construction	0	0	1	0
jordbävningen	the earthquake	0	0	1	0
jordbävningen	earthquake	0	0	1	0
melodier	melodies	0	0	1	0
byggd	built	0	0	1	1
demokratiska	democratic	0	0	1	0
bygga	building	0	0	1	0
bygga	build	0	0	1	1
indirekt	indirect	0	0	1	1
indirekt	indirectly	0	0	1	1
skadad	damaged	0	0	1	0
bara	only	0	0	1	1
skadan	damage	0	0	1	0
skadan	the damage	0	0	1	0
skadan	the hit	0	0	1	0
influerad	influenced	0	0	1	0
anderssons	anderssons	0	0	1	0
anderssons	andersson's	0	0	1	0
skadas	damaged	0	0	1	0
konstant	constant	0	0	1	1
folk	public	0	0	1	0
folk	people	0	0	1	1
influerat	influenced	0	0	1	0
dramatiskt	dramatic	0	0	1	0
dramatiskt	dramatically	0	0	1	1
assisterande	assistant	0	0	1	1
assisterande	assisted	0	0	1	0
assisterande	assisting	0	0	1	0
kris	crisis	0	0	1	1
nämner	mentions	0	0	1	0
nämner	names	0	0	1	0
skrivna	written	0	0	1	0
domkyrka	cathedral	0	0	1	1
domkyrka	abbey	0	0	1	0
krig	war	0	0	1	1
dramatiska	dramatic	0	0	1	0
dramatiska	dramatical	0	0	1	0
överlever	survives	0	0	1	0
sänktes	sunk	0	0	1	0
sänktes	reduced	0	0	1	0
koloni	colony	0	0	1	1
hårda	hard	0	0	1	0
hdmi	hdmi	0	0	1	0
producenten	the producer	0	0	1	0
producenten	producer	0	0	1	0
konto	account	0	0	1	1
konto	sign	0	0	1	0
turismen	tourism	0	0	1	0
turismen	the tourism	0	0	1	0
producenter	producers	0	0	1	0
diamanter	diamonds	0	0	1	0
filosofi	philosophy	0	0	1	1
astrid	astrid	0	0	1	0
tvingats	forced	0	0	1	0
tvingats	had	0	0	1	0
fauna	fauna	0	0	1	1
undre	lower	0	0	1	1
förstöra	destroy	0	0	1	1
förstöra	ruin; destroy	0	0	1	0
buddhistiska	buddhistic	0	0	1	0
buddhistiska	buddhist	0	0	1	0
ukraina	ukraine	0	0	1	0
metro	metro	0	0	1	1
innehar	holds	0	0	1	0
innehar	holding	0	0	1	0
innehas	held	0	0	1	0
innehas	occupied	0	0	1	0
innehav	possession	0	0	1	0
innehav	holdings	0	0	1	0
innehav	owning	0	0	1	0
anpassat	adapted	0	0	1	0
plattan	plate	0	0	1	0
plattan	the plate	0	0	1	0
inträffar	occur	0	0	1	0
inträffar	occurs	0	0	1	0
klädd	clothed	0	0	1	0
klädd	coated	0	0	1	0
inträffat	occurred	0	0	1	0
zlatan	zlatan	0	0	1	0
reda	find out	0	0	1	0
reda	find our	0	0	1	0
reda	out	0	0	1	0
gemenskap	fellowship	0	0	1	1
gemenskap	community	0	0	1	1
kristina	kristina	0	0	1	0
motor	engine	0	0	1	1
juryns	the jury's	0	0	1	0
juryns	jury	0	0	1	0
redo	ready	0	0	1	1
redo	prepared	0	0	1	0
lämnas	left	0	0	1	0
from	from	0	0	1	0
usa	the usa	0	0	1	0
usa	united states of america	0	0	1	0
usa	usa	0	0	1	0
fel	faults	0	0	1	0
fel	errors	0	0	1	0
fel	error	0	0	1	1
fem	five	0	0	1	1
hårdare	harder	0	0	1	1
hårdare	more severely	0	0	1	0
hårdare	tougher	0	0	1	0
vikingar	vikings	0	0	1	0
medicinskt	medical	0	0	1	0
utomstående	outside people; outsiders	0	0	1	0
utomstående	outside	0	0	1	0
utomstående	outsider	0	0	1	1
inlandet	inland	0	0	1	0
inlandet	the inland	0	0	1	0
sorg	grief	0	0	1	1
sorg	sad	0	0	1	0
andliga	spiritual	0	0	1	0
penis	penis	0	0	1	1
oerhört	tremendously	0	0	1	1
oerhört	extremely	0	0	1	0
hindrade	preventing	0	0	1	0
hindrade	prevented	0	0	1	0
nonsporting	non sporting	0	0	1	0
fungerar	functions	0	0	1	0
fungerar	works	0	0	1	0
slutade	quit	0	0	1	0
slutade	ending	0	0	1	0
beskriva	describe	0	0	1	1
automatiskt	automatic	0	0	1	0
black	black	0	0	1	0
monetära	monetary	0	0	1	0
beskrivs	described	0	0	1	0
flöde	feed	0	0	1	0
fälttåg	crusade	0	0	1	0
fälttåg	campaign	0	0	1	1
tar	takes	0	0	1	0
tas	is	0	0	1	0
tas	is taken	0	0	1	0
platser	points	0	0	1	0
platser	places	0	0	1	0
ställen	spots; places	0	0	1	0
ställen	places	0	0	1	0
ställen	stables	0	0	1	0
crick	cricket	0	0	1	0
crick	crick	0	0	1	0
engels	engels	0	0	1	0
ställer	running; causing	0	0	1	0
ställer	set	0	0	1	0
ställer	run (in election)	0	0	1	0
göta	göta	0	0	1	0
tag	while	0	0	1	0
hilton	hilton	0	0	1	0
stället	instead	0	0	1	0
stället	the place	0	0	1	0
tal	speech	0	0	1	1
kanadensiska	canadian	0	0	1	0
sir	sir	0	0	1	1
ondska	evil	0	0	1	1
utfärdade	issued	0	0	1	0
siv	siv	0	0	1	0
six	six	0	0	1	0
brian	brian	0	0	1	0
sig	to	0	0	1	0
sig	itself	0	0	1	1
öron	ear	0	0	1	0
öron	anxiety	0	0	1	0
öron	ears	0	0	1	0
sin	its	0	0	1	1
kostym	costume	0	0	1	1
kontroversiellt	controversial	0	0	1	0
företrädare	preferred traders	0	0	1	0
företrädare	representatives	0	0	1	0
roterande	rotating	0	0	1	1
framgångar	successes	0	0	1	0
framgångar	success	0	0	1	0
oavsett	whether	0	0	1	0
oavsett	regardless; whether; irrespective of	0	0	1	0
oavsett	regardless	0	0	1	1
tack	thanks	0	0	1	1
bertil	bertil	0	0	1	0
kategoriwikipediabasartiklar	category wikipedia basartiklar	0	0	1	0
kontroversiella	controversial	0	0	1	0
förbundskapten	manager	0	0	1	0
förbundskapten	coach	0	0	1	0
eritrea	eritrea	0	0	1	0
språkbruk	language (use); parlance; phraseology	0	0	1	0
språkbruk	parlance	0	0	1	1
språkbruk	language	0	0	1	0
light	light	0	0	1	0
självbiografi	autobiography	0	0	1	1
självbiografi	selfbiografi	0	0	1	0
sånger	songs	0	0	1	0
sången	the song	0	0	1	0
sången	song	0	0	1	0
centralorter	centers	0	0	1	0
centralorter	regional centers	0	0	1	0
kommunikationer	communications	0	0	1	0
jolie	jolie	0	0	1	0
jolie	jolies	0	0	1	0
besegrat	defeated	0	0	1	0
mekka	mecca	0	0	1	0
mekka	mecka	0	0	1	0
blandad	mixed	0	0	1	1
blandad	blended	0	0	1	0
skapande	building	0	0	1	0
skapande	creating	0	0	1	1
skapande	creative	0	0	1	1
elin	elin	0	0	1	0
elin	electrical	0	0	1	0
elit	elite	0	0	1	1
blandat	mixed	0	0	1	0
karlstad	karlstad	0	0	1	0
karlstad	phoenix	0	0	1	0
blandas	mixed	0	0	1	0
blandas	mixes	0	0	1	0
värld	world	0	0	1	1
spotify	spotify	0	0	1	0
stiga	rise	0	0	1	1
stiga	rising	0	0	1	0
terriers	terriers	0	0	1	0
invånarna	inhabitants	0	0	1	0
invånarna	inhabitatants; citizens'	0	0	1	0
invånarna	residents	0	0	1	0
befolkning	population	0	0	1	1
byn	village	0	0	1	0
permanent	permanent	0	0	1	1
märken	brands	0	0	1	0
märken	sign	0	0	1	0
genomsnittlig	average	0	0	1	1
datorn	the computer	0	0	1	0
datorn	pc	0	0	1	0
välmående	healthy	0	0	1	1
välmående	well-being; affluent	0	0	1	0
välmående	prosperous	0	0	1	1
carola	carola	0	0	1	0
cypern	cyprus	0	0	1	1
verkligen	real	0	0	1	0
verkligen	the reality	0	0	1	0
washington	washington	0	0	1	0
omedelbart	immediately	0	0	1	1
omedelbart	immediate	0	0	1	0
skickas	is sent	0	0	1	0
skickas	sent	0	0	1	0
skickas	any	0	0	1	0
skickar	sends	0	0	1	0
skickar	send	0	0	1	0
ön	island	0	0	1	0
ön	the island	0	0	1	0
satelliter	satellite	0	0	1	0
exempelvis	e.g.	0	0	1	0
brukar	usually	0	0	1	0
brukar	used to	0	0	1	0
komma	access	0	0	1	0
komma	get	0	0	1	0
billy	billy	0	0	1	0
uppvärmning	heating	0	0	1	1
uppvärmning	warming	0	0	1	0
förhåller	relate	0	0	1	0
förhåller	relationship	0	0	1	0
förhåller	relates	0	0	1	0
konungariket	kingdom	0	0	1	0
källorna	source	0	0	1	0
källorna	the sources	0	0	1	0
studios	studios	0	0	1	0
studios	the studio's	0	0	1	0
australiska	australian	0	0	1	0
färgade	colored	0	0	1	0
bröllopet	the wedding	0	0	1	0
bröllopet	wedding	0	0	1	0
barnets	the childs	0	0	1	0
barnets	the child's	0	0	1	0
barnets	child	0	0	1	0
kvarteret	quarter	0	0	1	0
kvarteret	the neighborhood	0	0	1	0
studion	studio	0	0	1	0
studion	the studio	0	0	1	0
kritik	criticism	0	0	1	1
kritik	critisism	0	0	1	0
kritik	critique; criticism	0	0	1	0
alger	algae	0	0	1	0
alger	algaes	0	0	1	0
blues	blues	0	0	1	0
uggla	owl	0	0	1	1
föreställning	performance	0	0	1	1
föreställning	present stall	0	0	1	0
minskad	decreased	0	0	1	0
minskad	reduced	0	0	1	0
längden	the length	0	0	1	0
längden	length	0	0	1	0
längden	lenght	0	0	1	0
hantverkare	craftsman	0	0	1	1
hantverkare	handy worker	0	0	1	0
fiktiva	fictitious	0	0	1	0
fiktiva	romantic	0	0	1	0
svar	answer	0	0	1	1
svar	response	0	0	1	1
waterloo	waterlo	0	0	1	0
waterloo	waterloo	0	0	1	0
består	consists of	0	0	1	0
består	beasts	0	0	1	0
består	exists	0	0	1	0
nobelpristagare	nobel laureate (-s); nobel prize winner (-s)	0	0	1	0
nobelpristagare	nobel laureates	0	0	1	0
minskat	decreased	0	0	1	0
minskat	reduced	0	0	1	0
minskat	has decreased	0	0	1	0
centralamerika	central america	0	0	1	0
minskar	diminishing	0	0	1	0
minskar	decrease	0	0	1	0
vulkanutbrott	volcanic eruption	0	0	1	0
vulkanutbrott	vulcano eruption	0	0	1	0
räddar	saves	0	0	1	0
räddar	saved	0	0	1	0
räddar	rescues	0	0	1	0
york	york	0	0	1	0
framgång	success	0	0	1	1
genomgår	undergoes	0	0	1	0
genomgår	undergoing	0	0	1	0
studioalbumet	studio album	0	0	1	0
philip	philip	0	0	1	0
ärkebiskopen	archbishop	0	0	1	0
domare	judge	0	0	1	1
fotbollslandslag	football team	0	0	1	0
fotbollslandslag	national football team	0	0	1	0
anslutning	connection	0	0	1	1
tyst	quiet	0	0	1	1
tyst	silent	0	0	1	1
varsin	(one) each	0	0	1	0
varsin	opposite	0	0	1	0
g	(g)	0	0	1	0
barns	childrens	0	0	1	0
barns	children	0	0	1	0
barns	child	0	0	1	0
via	via	0	0	1	1
via	through	0	0	1	0
framgår	will be seen	0	0	1	0
framgår	clear	0	0	1	0
framgår	is shown	0	0	1	0
adrian	adrian	0	0	1	0
familjens	the familys	0	0	1	0
familjens	family	0	0	1	0
tysk	german	0	0	1	1
rudolf	rudolph	0	0	1	0
rudolf	rudolf	0	0	1	0
revolutionens	revolution	0	0	1	0
revolutionens	the revolutions	0	0	1	0
isbn	isbn	0	0	1	0
brasilien	brazil	0	0	1	1
åkte	went	0	0	1	0
åkte	relegated	0	0	1	0
velat	wanted	0	0	1	0
kriterier	criteria	0	0	1	1
störningar	interruptions	0	0	1	0
störningar	disorder	0	0	1	0
störningar	disorders	0	0	1	0
ses	be	0	0	1	0
ses	are seen	0	0	1	0
påminner	reminds	0	0	1	0
påminner	out	0	0	1	0
bärande	wearing	0	0	1	0
bärande	leading	0	0	1	0
bärande	fundamental; wearing; supportive	0	0	1	0
regenter	monarchs	0	0	1	0
regenter	regents	0	0	1	0
skyddade	protected	0	0	1	0
enkelt	simple	0	0	1	0
enkelt	easy	0	0	1	1
övergick	transended	0	0	1	0
övergick	went over	0	0	1	0
övergick	switched	0	0	1	0
förväntade	expected	0	0	1	0
förmån	benefit	0	0	1	1
förmån	advantage; in favor of; benefit	0	0	1	0
meddelanden	messages	0	0	1	0
omfattning	extent	0	0	1	1
misslyckande	failure	0	0	1	1
innehålla	include	0	0	1	1
innehålla	contain	0	0	1	1
sankta	sankta	0	0	1	0
sankta	saint	0	0	1	1
diskutera	discussed	0	0	1	0
diskutera	discuss	0	0	1	1
mer	more	0	0	1	1
utsöndras	exudes	0	0	1	0
utsöndras	secrete	0	0	1	0
utsöndras	secreted	0	0	1	0
valda	chosen	0	0	1	0
övergå	transition	0	0	1	0
övergå	transend	0	0	1	0
vingar	wings	0	0	1	0
juli	july	0	0	1	1
vind	wind	0	0	1	1
stöds	supported	0	0	1	0
stöds	stood	0	0	1	0
stöds	is supported	0	0	1	0
resterande	remainder	0	0	1	0
resterande	remaining	0	0	1	1
franska	french	0	0	1	1
holland	holland	0	0	1	1
franske	the french	0	0	1	0
franske	french	0	0	1	0
birgitta	birgitta	0	0	1	0
tommy	tommy	0	0	1	0
algeriet	algeria	0	0	1	1
franskt	french	0	0	1	0
tomma	empty	0	0	1	0
kännetecken	characteristics	0	0	1	0
kännetecken	sign	0	0	1	0
kännetecken	distinction	0	0	1	0
tyskarna	the german	0	0	1	0
tyskarna	germans	0	0	1	0
tyskarna	the germans	0	0	1	0
händelse	suffix	0	0	1	0
händelse	handel	0	0	1	0
händelse	event	0	0	1	1
fyrtio	forty	0	0	1	1
bröderna	brothers	0	0	1	0
bröderna	the brothers	0	0	1	0
cohen	cohen - it's a name	0	0	1	0
cohen	cohen	0	0	1	0
störst	large	0	0	1	0
störst	most	0	0	1	0
benny	benny	0	0	1	0
ländernas	countries	0	0	1	0
ländernas	the countries	0	0	1	0
ländernas	countries'	0	0	1	0
blir	become	0	0	1	0
blir	is	0	0	1	0
farligt	dangerous	0	0	1	0
farligt	hazardly	0	0	1	1
ringen	ring	0	0	1	0
intervju	interview	0	0	1	1
storbritannien	great britain	0	0	1	1
storbritannien	uk	0	0	1	0
byggas	prevented	0	0	1	0
byggas	built	0	0	1	0
byggas	build	0	0	1	0
uppfann	invented	0	0	1	0
lopp	course	0	0	1	1
lopp	races	0	0	1	0
lopp	race	0	0	1	1
lopp	passage	0	0	1	1
besittning	dominion	0	0	1	1
besittning	possess	0	0	1	0
motorväg	autobahn	1	1	0	0
motorväg	motorway	1	1	0	1
motorväg	high way	1	0	1	0
motorväg	tyumen	1	0	1	0
motorväg	freeway	1	1	1	1
motorväg	tiumen	1	0	1	0
motorväg	highway	1	1	1	1
motorväg	interstate	1	1	0	0
kristi	kristi	0	0	1	0
kristi	christ	0	0	1	0
fördelningen	distribution	0	0	1	0
betydligt	considerably	0	0	1	1
betydligt	significant	0	0	1	0
förutsätter	assume	0	0	1	0
förutsätter	requires	0	0	1	0
förutsätter	assumes	0	0	1	0
centra	center	0	0	1	0
bära	carry	0	0	1	1
bära	mean	0	0	1	0
centre	center	0	0	1	0
centre	centre	0	0	1	0
who	who	0	0	1	0
landslaget	the national team	0	0	1	0
landslaget	team	0	0	1	0
intogs	was taken	0	0	1	0
intogs	was captured	0	0	1	0
staternas	states	0	0	1	0
staternas	the state's	0	0	1	0
bostäder	residences	0	0	1	0
bostäder	housing	0	0	1	0
förbi	past	0	0	1	1
förbi	past the	0	0	1	0
förbi	pass	0	0	1	0
regeringschef	head of government	0	0	1	1
regeringschef	government	0	0	1	0
miljontals	millions	0	0	1	0
enbart	only	0	0	1	0
judendomen	the judaism	0	0	1	0
judendomen	judaism	0	0	1	0
movie	movie	0	0	1	0
moberg	moberg	0	0	1	0
uefa	uefa	0	0	1	0
blandade	mixed	0	0	1	0
funktionella	functional	0	0	1	0
debatt	debate	0	0	1	1
planerna	the plans	0	0	1	0
planerna	plans	0	0	1	0
sämre	poor	0	0	1	0
sämre	samre	0	0	1	0
fann	found	0	0	1	0
julafton	chistmas eve	0	0	1	0
julafton	christmas eve	0	0	1	1
pastoral	pastoral	0	0	1	1
eiffeltornet	the eiffel tower	0	0	1	0
asterix	asterix	0	0	1	0
släkten	genera	0	0	1	0
släkten	the family	0	0	1	0
släkten	slaughter	0	0	1	0
filmer	films	0	0	1	0
filmer	movies	0	0	1	0
beroende	dependent	0	0	1	1
beroende	dependent on	0	0	1	0
beroende	depending	0	0	1	0
födelsedag	birthday	0	0	1	1
procent	percent	0	0	1	1
procent	per	0	0	1	0
heta	hot	0	0	1	0
heta	be named; be called	0	0	1	0
heta	be called	0	0	1	1
överlevt	survived	0	0	1	0
gudar	gods	0	0	1	0
hårdrocken	hard rock	0	0	1	0
presley	presley	0	0	1	0
hett	hot	0	0	1	0
överleva	survive	0	0	1	1
överleva	survival	0	0	1	0
överleva	over live	0	0	1	0
väldet	empire	0	0	1	0
väldet	violence	0	0	1	0
väldet	the rule	0	0	1	0
regler	rules	0	0	1	0
fötts	born	0	0	1	0
fötts	borned	0	0	1	0
samtycke	consent	0	0	1	1
samtycke	approval	0	0	1	0
tjänade	earning	0	0	1	0
tjänade	earned	0	0	1	0
dåtidens	past times	0	0	1	0
dåtidens	yesterdays	0	0	1	0
dåtidens	that time	0	0	1	0
förbjuda	forbid	0	0	1	1
förbjuda	ban	0	0	1	1
förbjuda	prohibiting	0	0	1	0
följdes	followed	0	0	1	0
följdes	was followed	0	0	1	0
strävhårig	hispid	0	0	1	0
strävhårig	wirehaired	0	0	1	0
utländsk	foreign	0	0	1	1
utländsk	foregin	0	0	1	0
uppgår	is	0	0	1	0
uppgår	shall amount	0	0	1	0
torka	dry	0	0	1	1
landets	the country's	0	0	1	0
landets	its	0	0	1	0
häcklöpning	hurdles	1	1	0	0
häcklöpning	hackopning	1	0	1	0
häcklöpning	hurdles race	1	0	1	0
häcklöpning	hurdling	1	1	0	0
häcklöpning	hurdle	1	0	1	1
häcklöpning	hacklopning	1	0	1	0
häcklöpning	coin	1	0	1	0
häcklöpning	hurdle race	1	1	0	0
häcklöpning	hurdle-race	1	0	1	1
mestadels	most of the time	0	0	1	0
mestadels	mostly	0	0	1	1
kvinnorna	the women	0	0	1	0
kvinnorna	women	0	0	1	0
färdas	travels	0	0	1	0
bäst	bast	0	0	1	0
bäst	best	0	0	1	1
nationernas	the nation's	0	0	1	0
nationernas	the nations	0	0	1	0
nationernas	nations	0	0	1	0
rikare	richer	0	0	1	0
lagerlöf	lagerlöf	0	0	1	0
lagerlöf	lagerlof	0	0	1	0
religiös	religious	0	0	1	1
theta	theta	0	0	1	0
funktion	function	0	0	1	1
upplysning	the enlightenment	0	0	1	0
upplysning	enlightenment	0	0	1	1
praktisk	practical	0	0	1	1
sydstaterna	the southern states	0	0	1	0
sydstaterna	southern states	0	0	1	0
sydstaterna	southern united states	0	0	1	0
menas	means	0	0	1	0
menas	mean	0	0	1	0
vandrar	wanders	0	0	1	0
vandrar	migrates	0	0	1	0
joe	joe	0	0	1	0
swift	swift	0	0	1	0
jon	jon	0	0	1	0
barrett	barett	0	0	1	0
barrett	barrett	0	0	1	0
grönt	green	0	0	1	1
allsvenskan	headlines	0	0	1	0
allsvenskan	allsvenskan	0	0	1	0
ingemar	ingemar	0	0	1	0
länders	countries	0	0	1	0
länders	countries'	0	0	1	0
länders	countrie's	0	0	1	0
teoretiker	say	0	0	1	0
teoretiker	theorists	0	0	1	0
infört	introduced	0	0	1	0
kolhydrater	carbons	0	0	1	0
kolhydrater	carbohydrates	0	0	1	0
april	april	0	0	1	1
brons	bronze	0	0	1	1
vattnets	water	0	0	1	0
vattnets	the water's	0	0	1	0
vattnets	the waters	0	0	1	0
bronx	bronx	0	0	1	0
bronx	the bronx	0	0	1	0
förmågan	the ability	0	0	1	0
släkt	pettigree	0	0	1	0
släkt	family	0	0	1	1
klasser	classes	0	0	1	0
betecknar	represent	0	0	1	0
betecknar	represents	0	0	1	0
betecknar	denotes	0	0	1	0
betecknas	denote	0	0	1	0
betecknas	labelled	0	0	1	0
betecknas	designate	0	0	1	0
kategorityska	category: german	0	0	1	0
demens	dementia	0	0	1	1
korruption	corruption	0	0	1	1
kämpa	fight	0	0	1	1
wall	wall	0	0	1	0
vittne	witness	0	0	1	1
publicerad	published	0	0	1	0
walt	walt	0	0	1	0
döptes	renamed; named	0	0	1	0
döptes	renamed	0	0	1	0
döptes	baptised	0	0	1	0
cirka	about	0	0	1	1
cirka	approximately	0	0	1	1
utsedd	appointed	0	0	1	0
styrkor	strenghts	0	0	1	0
styrkor	forces	0	0	1	0
publiceras	publishes	0	0	1	0
publiceras	will be published	0	0	1	0
publiceras	published	0	0	1	0
publicerat	published	0	0	1	0
själv	alone	0	0	1	0
själv	own	0	0	1	0
själv	himself	0	0	1	1
demografiska	demographic	0	0	1	0
demografiska	demographical	0	0	1	0
klara	clear	0	0	1	1
miljöer	environment	0	0	1	0
miljöer	environments	0	0	1	0
hindu	hindu	0	0	1	1
kopplade	connected	0	0	1	0
närma	move closer	0	0	1	0
närma	approach	0	0	1	0
närma	approximate	0	0	1	0
bbc	bbc	0	0	1	0
beskrivning	description	0	0	1	1
skånska	scanian dialect	0	0	1	0
skånska	scanian	0	0	1	0
skånska	skånska	0	0	1	0
klart	clear	0	0	1	1
klart	done	0	0	1	0
klart	finished	0	0	1	0
cry	cry	0	0	1	0
självmord	self-killing	0	0	1	0
självmord	suicide	0	0	1	1
strindbergs	strindberg's	0	0	1	0
strindbergs	strindberg	0	0	1	0
mike	micke	0	0	1	0
mike	mike	0	0	1	0
pengar	money	0	0	1	1
nickel	nickel	0	0	1	1
turneringen	the tournament	0	0	1	0
dominera	dominate	0	0	1	1
lutherska	lutheran	0	0	1	0
växt	plant	0	0	1	1
hms	hms	0	0	1	0
pjäsen	play	0	0	1	0
pjäsen	piece	0	0	1	0
neutrala	neutral	0	0	1	0
deklarerade	declared	0	0	1	0
plikter	duties	0	0	1	0
växa	growth	0	0	1	0
växa	grow	0	0	1	1
växa	wax	0	0	1	1
present	gift	0	0	1	1
släppte	released	0	0	1	0
problemen	problems	0	0	1	0
problemen	the problems	0	0	1	0
officiell	official	0	0	1	1
officiell	authentic	0	0	1	0
anpassa	adjust	0	0	1	1
anpassa	adapt	0	0	1	1
will	will	0	0	1	0
östman	Östman	0	0	1	0
yngre	younger	0	0	1	1
wild	wild	0	0	1	0
madeleine	madeleine	0	0	1	0
kommande	upcoming	0	0	1	0
sagan	story	0	0	1	0
uppfattning	view	0	0	1	0
uppfattning	understanding	0	0	1	1
ställe	stalle	0	0	1	0
ställe	place	0	0	1	1
tränga	push (aside)	0	0	1	0
tränga	cut in	0	0	1	0
tränga	permeate	0	0	1	0
gemensamt	single	0	0	1	0
gemensamt	in common	0	0	1	1
syftar	refers	0	0	1	0
syftar	seek to	0	0	1	0
syftar	refer	0	0	1	0
fötterna	feet	0	0	1	0
fötterna	their feet	0	0	1	0
fötterna	the feet	0	0	1	0
decennierna	decades	0	0	1	0
decennierna	the decades	0	0	1	0
motiv	subjects	0	0	1	0
motiv	motif	0	0	1	1
jehovas	jehovas	0	0	1	0
jehovas	jehova's	0	0	1	0
halt	content	0	0	1	1
halt	stop; level	0	0	1	0
halt	stop	0	0	1	0
ramels	ramel's	0	0	1	0
överlevnad	survival	0	0	1	0
varar	duration	0	0	1	0
varar	lasts	0	0	1	0
föda	feed	0	0	1	1
föda	give birth; food	0	0	1	0
föda	give birth	0	0	1	0
buddhism	buddhism	0	0	1	1
behövdes	required	0	0	1	0
pojkar	boys	0	0	1	0
samband	connection	0	0	1	1
inch	inches	0	0	1	0
skickade	sent	0	0	1	0
gett	given	0	0	1	0
gett	gave	0	0	1	0
annekterade	annexed	0	0	1	0
annekterade	annexation	0	0	1	0
tvister	conflicts	0	0	1	0
tvister	disputes	0	0	1	0
mottagande	host	0	0	1	0
mottagande	reception	0	0	1	1
vänder	turn	0	0	1	0
vänder	vander	0	0	1	0
vänder	face	0	0	1	0
romeo	romeo	0	0	1	0
konst	art	0	0	1	1
konst	srt	0	0	1	0
romer	romani people	0	0	1	0
romer	roma	0	0	1	0
student	student	0	0	1	1
raka	straight	0	0	1	0
översättningar	translations	0	0	1	0
misstag	mistake	0	0	1	1
misstag	error	0	0	1	1
klubbar	clubs	0	0	1	0
vilar	rests	0	0	1	0
banden	bands	0	0	1	0
banden	bander	0	0	1	0
banden	the bound	0	0	1	0
färgen	color	0	0	1	0
färgen	the color	0	0	1	0
ekosystem	ecosystem	0	0	1	1
ekosystem	eco system	0	0	1	0
individens	individual's	0	0	1	0
individens	the individual's	0	0	1	0
färger	color	0	0	1	0
färger	farger	0	0	1	0
färger	colors	0	0	1	0
english	english	0	0	1	0
bandet	band	0	0	1	0
organisationens	organization	0	0	1	0
organisationens	the organizations	0	0	1	0
biologisk	biological	0	0	1	1
singeln	single	0	0	1	0
singeln	singeln	0	0	1	0
mfl	etc	0	0	1	0
mfl	etc.	0	0	1	0
uppkommer	arises	0	0	1	0
uppkommer	resulting	0	0	1	0
uppkommer	arises; generated	0	0	1	0
känner	kanner	0	0	1	0
känner	knows	0	0	1	0
känner	know	0	0	1	0
rachels	rachels	0	0	1	0
rachels	rachel's	0	0	1	0
erfarenheter	experiences	0	0	1	0
erfarenheter	experience	0	0	1	0
patrik	patrik	0	0	1	0
antisemitism	antisemitism	0	0	1	1
rocken	the rock	0	0	1	0
rocken	rock	0	0	1	0
brutit	cut; break	0	0	1	0
brutit	broken	0	0	1	0
mytologiska	mytholigical	0	0	1	0
mytologiska	mythological	0	0	1	0
ändrar	changing	0	0	1	0
ändrar	changes	0	0	1	0
ändrar	change	0	0	1	0
jarl	earl	0	0	1	0
jarl	jarl	0	0	1	1
genombrottet	break-through	0	0	1	0
genombrottet	breakthrough	0	0	1	0
alldeles	completely	0	0	1	1
alldeles	altogether	0	0	1	1
hoppa	skip	0	0	1	1
hoppa	drop out	0	0	1	0
sky	sky	0	0	1	1
engelsk	english	0	0	1	1
ske	be	0	0	1	0
ske	happen	0	0	1	1
resultat	results	0	0	1	1
resultat	result	0	0	1	1
fyller	turns	0	0	1	0
fyller	play	0	0	1	0
fyller	turn; fill	0	0	1	0
sanskrit	sanskrit	0	0	1	1
stolpiller	web	1	0	1	0
stolpiller	network	1	0	1	0
stolpiller	suppositary	1	0	1	0
stolpiller	pauropoda	1	0	1	0
stolpiller	suppository	1	1	0	1
stolpiller	suppositories	1	1	0	0
stolpiller	stolpills	1	1	0	0
hotade	threatened	0	0	1	0
psykoser	psychoses	0	0	1	0
psykoser	psychosis	0	0	1	0
jordbävning	earthquake	0	0	1	1
agerande	acting	0	0	1	0
agerande	behavior	0	0	1	0
landshövding	county governor	0	0	1	0
landshövding	govenror	0	0	1	0
landshövding	governor	0	0	1	1
förekomsten	existence	0	0	1	0
förekomsten	presence	0	0	1	0
know	know	0	0	1	0
press	press	0	0	1	1
psykosen	psychosis	0	0	1	0
psykosen	the psychosis	0	0	1	0
institut	institute	0	0	1	1
institut	institution	0	0	1	1
georges	georges	0	0	1	0
budet	the bid	0	0	1	0
budet	the commandment	0	0	1	0
miami	miami	0	0	1	0
djupa	deep	0	0	1	0
huruvida	whether	0	0	1	1
gorbatjov	gorbachev	0	0	1	0
gorbatjov	gotbatjov	0	0	1	0
finansieras	financed	0	0	1	0
finansieras	funded	0	0	1	0
finansieras	finansed	0	0	1	0
djupt	deeply	0	0	1	1
djupt	deep	0	0	1	1
serbiska	serbian	0	0	1	0
säkerheten	the security	0	0	1	0
säkerheten	safety	0	0	1	0
tjeckoslovakien	czechoslovakia	0	0	1	0
handeln	trade; commerce	0	0	1	0
handeln	trade	0	0	1	0
bibliska	biblican	0	0	1	0
bibliska	biblical	0	0	1	0
aktier	share	0	0	1	0
aktier	stock	0	0	1	0
handels	commercial	0	0	1	0
handels	trade	0	0	1	0
förorter	suburbs	0	0	1	0
självstyre	autonomy	0	0	1	0
självstyre	self-governance	0	0	1	0
självstyre	self-government	0	0	1	0
star	star	0	0	1	0
empire	empire	0	0	1	0
skandinavien	scandinavia	0	0	1	1
genomsnitt	average	0	0	1	1
planering	planning	0	0	1	1
trianglar	with triangles	0	0	1	0
trianglar	traingles	0	0	1	0
gammalt	old	0	0	1	0
tvfilm	tv-movie	0	0	1	0
tvfilm	tv film	0	0	1	0
tvfilm	tv movie	0	0	1	0
undviker	avoids	0	0	1	0
undviker	avoid	0	0	1	0
björn	bear	0	0	1	1
björn	björn	0	0	1	0
setts	observed	0	0	1	0
setts	seen	0	0	1	0
mankell	mankell	0	0	1	0
spår	track	0	0	1	1
spår	pairs	0	0	1	0
stieg	stieg	0	0	1	0
förbindelser	connections	0	0	1	0
förbindelser	relations	0	0	1	0
sjunker	flag	0	0	1	0
sjunker	sinks	0	0	1	0
markera	mark	0	0	1	1
efteråt	afterwards	0	0	1	1
decennium	decade	0	0	1	1
mitt	my	0	0	1	1
mitt	center	0	0	1	1
omskärelse	circumcision	0	0	1	1
slut	end	0	0	1	1
slut	out	0	0	1	1
sommarspelen	summer games	0	0	1	0
sommarspelen	summer olympics	0	0	1	0
eran	era	0	0	1	0
lämnar	leaves	0	0	1	0
ljung	heather	0	0	1	1
lämnat	left	0	0	1	0
pressfrihetsindex	press freedom index	0	0	1	0
pressfrihetsindex	pressfrihetsindex	0	0	1	0
substantiv	noun	0	0	1	1
or	or	0	0	1	0
oberoende	independent	0	0	1	1
avsnittet	section	0	0	1	0
avsnittet	episode	0	0	1	0
spektrum	spectra	0	0	1	0
spektrum	spectrum	0	0	1	1
saken	the thing	0	0	1	0
saken	matter	0	0	1	0
saken	the matter	0	0	1	0
saker	things	0	0	1	0
saker	items	0	0	1	0
avsnitten	the episodes	0	0	1	0
avsnitten	sections	0	0	1	0
avsnitten	chapters	0	0	1	0
own	egen	0	0	1	0
sjöfart	sea voyage	0	0	1	0
sjöfart	navigation	0	0	1	1
sjöfart	maritime	0	0	1	0
egna	own	0	0	1	0
egna	custom	0	0	1	0
floder	rivers	0	0	1	0
stanna	stop	0	0	1	1
stanna	stay	0	0	1	1
öl	beer	0	0	1	1
tillbringade	spent	0	0	1	0
mälaren	mälaren	0	0	1	0
sektorn	sector	0	0	1	0
sektorn	the sector	0	0	1	0
floden	river	0	0	1	0
floden	the river	0	0	1	0
vidta	take	0	0	1	1
hänvisa	reference	0	0	1	0
hänvisa	refer	0	0	1	1
flyger	flies	0	0	1	0
flyger	flying	0	0	1	0
hänt	suspension	0	0	1	0
hänt	happened	0	0	1	0
glukos	glucose	0	0	1	1
folkpartiet	peoples party	0	0	1	0
folkpartiet	liberal party	0	0	1	0
konstruktion	construction	0	0	1	1
konstruktion	structure	0	0	1	0
van	van	0	0	1	0
val	elections	0	0	1	0
val	election	0	0	1	1
val	choice	0	0	1	1
försvarets	defense	0	0	1	0
försvarets	forsvarets	0	0	1	0
försvarets	the defence's	0	0	1	0
missionärer	missioners	0	0	1	0
missionärer	missioner	0	0	1	0
missionärer	missionaries	0	0	1	0
vad	as	0	0	1	0
vad	what	0	0	1	1
smeknamnet	nickname	0	0	1	0
värmlands	värmlands	0	0	1	0
värmlands	varmlands	0	0	1	0
värmlands	hot countries	0	0	1	0
valuta	currency	0	0	1	1
valuta	exchange	0	0	1	0
var	was	0	0	1	0
regisserad	directed	0	0	1	0
regisserad	produced	0	0	1	0
bevarade	preserved	0	0	1	0
nordamerikanska	north american	0	0	1	0
lundell	lundell	0	0	1	0
identifierade	identified	0	0	1	0
förmedla	pass; express; mediate	0	0	1	0
förmedla	pass	0	0	1	0
granne	neighbour	0	0	1	1
granne	neighbor	0	0	1	1
förekom	ods	0	0	1	0
förekom	was	0	0	1	0
hänger	depends	0	0	1	0
hänger	hanger	0	0	1	0
öken	ok	0	0	1	0
öken	desert	0	0	1	1
hundratal	100	0	0	1	0
hundratal	hundred	0	0	1	0
krigsslutet	end of war; war's end	0	0	1	0
krigsslutet	end of the war	0	0	1	0
tänker	thinking	0	0	1	0
tänker	tankers	0	0	1	0
karta	map	0	0	1	1
karta	maps	0	0	1	0
made	made	0	0	1	0
erkänner	admits	0	0	1	0
erkänner	recognize	0	0	1	0
följs	followed	0	0	1	0
rybak	rybak	0	0	1	0
uppfattningar	opinions	0	0	1	0
uppfattningar	perceptions	0	0	1	0
arne	arne	0	0	1	0
tema	theme	0	0	1	1
följa	following	0	0	1	0
följa	follow	0	0	1	1
filip	filip	0	0	1	0
filip	phillipe	0	0	1	0
följd	following	0	0	1	0
följd	consequence	0	0	1	1
följd	effect	0	0	1	0
inledning	introduction	0	0	1	1
inledning	the beginning	0	0	1	0
kuriosa	bric-a-brac	0	0	1	0
kuriosa	curiosities	0	0	1	0
kuriosa	trivia	0	0	1	0
reaktorn	the reactor	0	0	1	0
reaktorn	reactor	0	0	1	0
problemet	problem	0	0	1	0
problemet	the problem	0	0	1	0
stormakter	world powers	0	0	1	0
stormakter	great power	0	0	1	0
stormakter	superpowers	0	0	1	0
kroatiska	croatian	0	0	1	0
pjäser	plays	0	0	1	0
pjäser	checkers	0	0	1	0
söderut	further south	0	0	1	0
söderut	south	0	0	1	0
låter	let	0	0	1	0
runor	runes	0	0	1	0
kant	kant	0	0	1	0
kant	edge	0	0	1	1
fullständigt	completely	0	0	1	1
fullständigt	full	0	0	1	1
illinois	illinois	0	0	1	0
rike	kingdom	0	0	1	1
book	book	0	0	1	0
normal	normal	0	0	1	1
porträtt	portraits	0	0	1	0
porträtt	portrait	0	0	1	1
fullständiga	full	0	0	1	0
fullständiga	complete	0	0	1	0
äldre	old	0	0	1	0
äldre	older	0	0	1	1
ursprunget	origin	0	0	1	0
ursprunget	the origin	0	0	1	0
intresse	interest	0	0	1	1
juni	june	0	0	1	1
tolkas	is interpreted	0	0	1	0
tolkas	interpretation	0	0	1	0
tolkas	interpret	0	0	1	0
tolkar	interprets	0	0	1	0
tolkar	views	0	0	1	0
shakespeares	shakespeare's	0	0	1	0
shakespeares	shakespeare	0	0	1	0
risker	risk	0	0	1	0
risker	risker	0	0	1	0
risker	risks	0	0	1	0
personligen	individual	0	0	1	0
personligen	personally	0	0	1	1
taube	taube	0	0	1	0
margaret	margaret	0	0	1	0
förmodligen	probably	0	0	1	0
förmodligen	presumably	0	0	1	1
markant	considerably	0	0	1	0
markant	markedly	0	0	1	0
markant	marked	0	0	1	1
risken	the risk	0	0	1	0
risken	risk	0	0	1	0
fransmännen	the french	0	0	1	0
fransmännen	frenchman	0	0	1	0
fransmännen	french	0	0	1	0
cliff	cliff	0	0	1	0
stadens	the town's	0	0	1	0
stadens	the citys	0	0	1	0
stadens	city's	0	0	1	0
knappast	hardly	0	0	1	1
knappast	dead	0	0	1	0
spontant	spontaneous	0	0	1	0
spontant	spontaneously	0	0	1	0
bysantinska	byzantine	0	0	1	0
blogg	blog	0	0	1	0
tidning	newspaper	0	0	1	1
tidning	journal	0	0	1	1
