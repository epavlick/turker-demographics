vanligast	most,most usual,most common,
nordisk	norse,nordic,
uppemot	up,
stammarna	tribes,strains,
arternas	the species,
jihad	johad,jihad,
invandrare	immigrants,
albumet	album,
slå	hit,sla,
lord	lord,
effektivt	effective,
lyckats	succeeded,
organisation	body,organization,
regional	regional,
upptar	occupies,
lämnades	was,
portugals	portugal,
dels	both,partly,
skicklig	proficient,
medelhavet	mediterranean,
helsingborg	helsingborg,
haber	haber,
befogenheter	authorities,
triangelns	triangle,
urskilja	distinguish,
sovjetisk	soviet,sovjetic,sovietic,
miller	miller,
sture	sture,
sammansatta	composed,
selassie	selassie,
ungerns	hungary,
upprätthåller	maintains,maintaining,
åsikten	the opinion,view,
breddgraden	latitude,
fossil	fossil,
punkt	point,
jönsson	jönsson,
filosofer	philosopher,
aten	athens,
hårda	hard,
vägrar	refuses,
filosofen	the philosopher,
motståndsrörelsen	resistance,
regnskog	rain forest,rainforest,
herr	mr,
föräldrarna	the parents,parents,
valrörelsen	election campaign,the election campaign,
bipolär	bipolar,
kids	kids,
demokratier	democracies,
vicepresident	vice president,
finska	finnish,
robin	robin,
miljarder	billions,
karin	karin,
tillverkningen	production,
systematiska	systematic,
unik	unique,
norsk	norwegian,
välkänd	well known,
systematiskt	systematic,
ansluta	join,connect,
dna	dna,
sjukdomen	disease,
strikt	strict,
fuktiga	futiga,
betraktats	considered,been seen,(been) viewed,
dns	dns,
fuktigt	moist,
musik	music,
befolkningstillväxten	population growth,the population growth,the growth of population,
holm	holm,
politiker	politicians,
slutligen	back end,
temperaturen	temperature,
kalksten	limestone,
temperaturer	temperature,
ofta	usually,often,
avancerad	advanced,
styrkan	strength; unit; force,strength,
köpa	buy,purchasing,
befolkningsutveckling	population development,population growth,
stommen	body,
syrgas	oxygen,
kapitalismen	capitalism,
vänner	friendas,friends,
igelkottar	hedgehogs,
kallare	colder,
hov	court,
how	how,
hot	hot,
hos	of,in; with,
folkmusik	folk music,
typen	type,
fylla	fill,
inrikes	domestic,
trettioåriga	13 year olds,thirty year's (war),
pengar	money,
barbro	barbro,
fyllt	filled,
objekt	objects,object,
turkiet	turklet,turkey,
sankt	st.,
typer	characters,types,
stormaktstiden	great power period,
isär	ice,apart,
deutsche	deutsche,
vart	each,
varv	shipbuilding,
ormar	snakes,
dalí	dali,
organismen	the organism,
vare	either,
varg	wolf,
organismer	organism,organisms,
vara	be,
omvandlas	convert,converted,
mabel	mabel,
befälhavare	commander,
publicerade	published,
besläktade	related,
nutida	present(-day); contemporary,present,
wales	wales,
målade	painted,
assyriska	assyrian,
fil	file,
avgå	resign,
väte	hydrogen,
hemlighet	secretly,
säljande	selling,
bestämmer	decide,
hänga	hang,
närliggande	adjacent,
utvecklat	developed,
utlänningar	foreigners,
utvecklar	develops,development speaker,
framsteg	progress,
terrorister	terrorists,
tingslag	things type,
debut	debut,
tillgängligt	available,
andrew	andrew,
ingrid	ingrid,
tillgängliga	available,
uppnådde	met,achieved,
talade	spoken,spoke,
angola	angola,
serier	comics,
allan	allan,
utvecklandet	development,
serien	the series,
velat	wanted,
axelmakterna	the axis,axis,
varken	either,
slovenien	slovenia,
tornet	tower,the tower,
debatter	debates,
anarkister	anarchists,
metallica	metallica,
arbetsplats	workplace,
ägnade	dedicated,
sannolikt	probably,probable,
sysselsätter	employs,
okända	unknown,
malmös	malmö's,malmö,
sydost	south east,
givetvis	naturally,
avsett	regard,
övre	upper,
avlägsna	remove,
förespråkar	occurring crackles,advocates,
vågade	dared,
ära	honor,
bitter	bitter,
förändringarna	changes,change,
senaten	senate,
bokstäverna	the letters,letters,
placerade	put,placed (in),
nirvana	nirvana,
påverkad	influenced,affected,
ahmed	ahmed,
skatter	taxes,
upphov	origin,source,
tyckte	find,
sköt	forwarder,shot,
tree	tree,
förstaplatsen	first place,
sorters	kinds of,kinds,
påverkat	influenced,affected,
varje	each,
påverkar	affecting,
påverkas	affected,
obligatorisk	obligatory,
hud	skin,
försörja	support,
assistent	assistant,
kriterierna	criteria,
boston	boston,
dricker	drinking,drink,
filosofisk	philosophical,philosophic,
halva	half,
joakim	joakim,
trakten	the region,region,
fasta	solid,
kroatien	croatia,
krigsmakt	military power,armed forces,
skaffa	obtain,
förhärskande	dominant,
hjälpmedel	resources,means agent,
katalonien	catalonia,
victoria	victoria,
gallagher	gallagher,
medlemsstaterna	member states,
anteckningar	notes,
bedriva	carry,
eftersom	because,
thriller	thriller,
övertog	took over,
annars	else,
singer	singer,
morgon	tomorrow,morning,
öland	oland,
camp	camp,
utmärkande	characteristic,distinguishing,
förlorar	loss,loses,
översatt	translated,
förlorat	lost,
producent	producer,
passerade	passed,
singel	single,
ned	bottom,
majs	corn,
ungar	babies,kids; offsprings; young,
representanter	representatives,
anorektiker	anorectic,
bandmedlemmar	band members,
nacka	nacka,
pris	price,
madeira	madeira,
teater	theatre; theater,theater,
louise	louis,louise,
populärkultur	popular culture,pop-culture,
buss	bus,
than	than,
övergår	surpasses,exceed,
rico	rico,
bush	bush,
rice	rice,
mottog	received,
lastbilar	trucks,
storbritanniens	united kingdom,uk,
årsdag	anniversary,
metoder	methods,
upprätta	up,
dansk	danish,
bensin	gasoline,
lyssna	listening,
balans	balance,
innebörd	meaning,
hantverk	crafts,
kallt	cold,coldly,
utgåvan	edition,the edition,
uppgift	data,
framfördes	framfordes,were,
genomsnittet	average,the average,
release	release,
kalla	cold,
ovtjarka	ovtjarka,
blev	became,
flagga	flag,
skulle	could,would,
skriva	write,
bygger	based,(is) building (on),
arlanda	arlanda,
skrivs	written,
nuförtiden	nowadays,
hedersdoktor	honorary doctor,
manson	manson,
förhindra	prevent,
upphovsrätt	copyright,
sundsvalls	sundsvall,(city of) sundsvall's,
figur	figure,
sista	last,
siste	last,
österrike	austria,
ringa	call,
rollen	the role,
henrik	henrik,
ställning	position,stall,
lanserades	launched,was launched,
konsekvens	impact,
tilldelades	awarded,
öst	east,
centralort	central city,regional centre,
tillämpas	applied,
huvudet	head,
country	country,
sparta	spartans,sparta,
följas	followed,
pitt	pitt,
edgar	edgar,
nederlag	defeat,
nordiskt	nordic,
genus	genus,
logik	logic,
aktuell	current,
igelkotten	the hedgehog,
folkmordet	genocide,
uttal	pronunciation,
baháulláh	bahaullah,
ana	ana,
fra	fra,
union	union,
avgörande	settling,decisive,essential,
fri	free,
operationer	operations,
socialistiskt	socialist,
årtionde	decade,
fru	madam,mrs.,
arbetslösheten	unemployment,
verktyg	tool,tools,
barndom	childhood,
life	life,
café	coffeehouse,café,
snittet	average,the average,
huvudstäder	capital cities,capitals,
ändrade	changed,modified,
arkiv	archives,
närvarande	present,
dave	dave,
chile	chile,
övergripande	over arching,overall,general,
chili	chili,
parterna	parties,
intag	intake,
uttryck	expression,
frankrikes	france's,
castro	castro,
klarade	passed,
organisera	organizing,
kontraktet	the contract,
tintin	tintin,
åke	åke,
brister	failures,
gärna	i'd love to,
desto	the,ever,
stämma	meeting,
player	player,
tänkare	thinker,
bristen	lack of,
madonna	madonna,
tät	compact,sealed,
memorial	memorial,
serbisk	serbian,
tillhandahåller	provides,
vrida	twist,turn,turning,
foton	images,photos,
omkring	about,
european	european,
kina	china,
materiell	material,
funktionen	the function,
topp	top,
värde	value,
tunn	thin,
föras	taken to,
synder	sins,
tung	heavy,
zeeland	zealand,
centraleuropa	central europe,
grundlag	constitution,
manteln	the mantle,mantle,
köra	drive,
koloniseringen	the colonization,colonization,
capitol	capitol,
dödsoffer	casualty,death victim,victim,
biskop	bishop,
krigsmakten	armed forces,
körs	running,being driven,
birmingham	birmingham,
utrotning	extinction,
döda	dead,
givit	gave,
matteus	matteus,
han	he,
grafit	graphite,
vetenskapsmän	scientist,scientists,
bnp	gnp,
muhammeds	mohammed's,muhammad,muhammed's,
huvud	head,main,
hette	named,hatte,
har	has,have,
hat	hatred,
hav	sea,
inne	inside,in,
underliggande	underlying,
ovanpå	top,
svensson	svensson,
narkotika	drug,narcotics,
livsstil	life style,lifestyle,
dagar	says,day,
melodifestivalen	eurovision song contest,
uppmärksammade	observed,noted,noticed,
bobby	bobby,
sedlar	bills,
alice	alice,
konsert	concert,
residensstad	city of residence,county seat,
sebastian	sebastian,
ola	ola,
people	people,
reagera	reacting,reaching,
islamisk	islamic,
parlamentarisk	parliamentary,
delade	divided,
fot	ft,
varierande	varied,
angränsande	adjacent,
utser	chooses,appoints,
utses	is appointed,
akademi	academy,
litterära	literary,
myndigheter	agencies,
annan	another,
neptunus	neptunes,
stefan	stefan,
påminner	out,
binder	tie,
olympiska	olympic,
möjligheterna	possibilities,the possibilities,
myndigheten	the authority,
annat	other; another,
army	army,
o	oh,
mynnar	opening,
klubben	club,
stjärna	star,
nixon	nixon,
tillverkare	producer,
hänt	happened,
delvis	partial,
döpte	baptized,
marshall	marshall,
ström	stream,
lagliga	legal,
son	son,
psykiskt	psychic,mentally,
delarna	the parts,parts,
america	america,
artikeln	the article,
hantera	handle,
nova	nova,
joseph	joseph,
jane	jane,
happy	happy,
saltkråkan	salt crow,saltkrakan,
jönköpings	jönköpings,jonkopings,
förhållandet	the ratio,relationship,
förhållanden	relationships,
öppet	open,
verde	verde,
tigern	tiger,
förväntningar	expectations,
drabbat	affected,
drabbas	suffer,troubled with,
polska	polish,
pest	plague,
syftet	purpose,
fansen	fans,
moderna	modern,
föregångare	predecessor,
konung	king,
lunds	lund's,lund,
låtar	songs,
modernt	modern,
krävde	demanded,
ericsson	ericsson,
astronomiska	astronomical,
huvudperson	main character,
dotter	daughter,
protester	protests,
republik	republic,
roll	role,
olja	oil,
reggae	reggae,
avskaffades	was abolished,abolished,
bostadsområden	residential areas,
palme	palme,
blått	blue,
vintrarna	winters,
modell	model,
utbildade	educated,formed,
danske	danish,dane,
tävling	competition,
danska	danish,
sällan	rare,
laddade	charged,
perioden	period,time,
kategorifödda	category born,category: born,
förtjust	fond,
tänderna	teeth,
herren	the lord,
perioder	period,periods,
erkända	acknowledged,recognized,
skatt	tax,
erkände	confession,acknowledged,
oss	us,
ost	cheese,
uppgifter	tasks,data,
stödjer	support,
avalanche	avalanche,
uppgiften	task,
atombomben	atomic bomb,
stålgemenskapen	steel community,
inkomst	income,
behåller	keeps,
fängelset	prison,
intresserade	interested,
vem	who,
framställa	produce,the installation,
bosnien	bosnia,
individer	individuals,
choice	choice,
individen	individual,
framställs	is depicted,prepared,
skillnaderna	the differences,differences,
kusterna	the coasts,coasts,
initiativ	initiative,
lägre	lower,
inhemska	native,
myntade	coined,
saab	saab,
oppositionen	opposition,
team	team,
uppskattningsvis	estimated,
årig	minor,
jämnt	even,
nybildade	newly formed,newly established,
scen	scene,
jämna	even,
firandet	the celebration,
måne	moon,
elton	elton,
köp	purchase,
kör	run,
kunskapen	knowledge,
beskydd	conservation,protection,
axel	axel,
bosatte	settled,
kön	gender,
kusten	the coast,coast,
katter	cats,cat,
berättelsen	story,the story,
provinserna	provinces,the provinces,
galileo	galileo,
skydd	protection,
budskapet	message,the message,
katten	the cat,
huvudsakliga	main,
studien	study,the study,
genomgående	consistently,pervading,
hälft	half,
landslag	national team,
studiet	the study,
studier	studies,
publicera	publish,
presenterade	presented,
smitta	infection,
samlar	salmar,
samlas	together,
änglar	angels,
vuxna	adult,
emellan	inbetween; between,between,
judarna	the jews, therefore,
positivt	positive,
samlag	intercourse,
effektiv	effective,
ställt	taken,set,
ställs	is,stalls,
dagars	day's,day,days,
hår	hair,
tillträdde	assumed,took,tilltradde,
ställe	stalle,place,
hål	hole,hal,
tabellen	the chart,
grönt	green,
straffet	penalty,the punishment,
kunskap	knowledge,
gröna	green,
phoebe	phoebe,
påvisa	detection,show,prove,
locka	attract,tempt,
missförstånd	misunderstandings,
locke	locke,
släktskap	relationship,kinship,
inkluderade	included,
rädda	save,lot of,
porträtt	portraits,portrait,
utnyttjade	utilized,used,
korta	short,
milda	mild,
årligen	annually,yearly,annual,
skikt	layer,
svenskan	swedish,the swede,
storleken	size,
trigonometriska	trigonometric,
levande	live,
riksdagen	the parliament,
gigantiska	gigantic,
kungens	king,the king's,
löpande	assembly,conveyor (belt),
ipredlagen	ipred act,
nyligen	recently,
data	data,
epost	e-mail,email,
stress	stress,
natural	natural,
bergarter	rocks,
undervisning	undervising,education,
påstod	claimed,said,
ss	ss,
sv	sw,south west,
sk	so called,
so	so,
vika	fold,
se	see,
resulterar	results,
vintrar	winters,
resulterat	resulted in,
professorn	the professor,
kong	(hong) kong,
antingen	presumably,either,
torg	square,
ingvar	ingvar,
utsätts	exposed,
jim	jim,
turnera	tour,
ersätts	replaced,
faderns	his father,
monopol	monopoly,
personlig	personal,
britter	britons,
pågick	lasted,
änden	end,spirit,
äldste	elders,eldest,
musiken	the music,music,
äldsta	oldest,
matcher	matches,games,
nation	nation,
matchen	the game,
kategoripersoner	category of persons,
efterföljande	subsequent,
twilight	twilight,
musiker	musicians,
atmosfär	atmospheric,
lockar	attracts,curls,
förväxlas	mixed up (with),confused,mistaken,
sidor	pages,sides,
säga	say,
tränade	trained,
dominerar	dominate,
domineras	dominated,
runstenar	runestones,rune stones,
sägs	said (to be),
dominerat	dominated,
födelsedag	birthday,
prisma	prism,
dynamiska	dynamic,
greker	greeks,
står	standing,
förstöra	destroy,ruin; destroy,
stål	steel,rate,
hinduer	hindus,
krav	requirement,conditions,
kött	cones,meat,
riktigt	real,right,
ockupationen	occupation,
sjuka	disease,
orsakar	causes,
riktiga	real,
bränder	fires,
internet	internet,
roterar	rotates,
bla	blah,among others,
sfären	spheres,
garantera	ensure,guarantee,
vård	vard,nursing,healthcare,
våra	our,
singlar	singles,
sålde	sold,sells drinks,
bytt	changed,switched,
byts	changed,replaced,
sålda	sold,salda,
väster	west,
vårt	each,
kolonier	colonies,
dramaten	dramaten,
byte	change of,bytes,
byta	switch,change,trade,
föreställning	performance,
pund	pound,
artister	performers,artists,
punk	punk rock,punk,para,
flandern	flanders,
solna	solna,
artisten	the artist,artist,
gordon	gordon,
främst	foremost; primarily; chiefly,all,
givits	given,
förmån	benefit,advantage; in favor of; benefit,
hård	hard,
potter	potter,
beethoven	beethoven,
tsunamier	tsunamis,
open	open,
ont	bad,
urin	urine,
city	city,
flytande	floating,liquid,
teologi	theology,
skådespelarna	actors,
råolja	crude oil,
intill	adjacent to,adjacent,
sjö	naval,
nästa	next,
williams	williams,
animerade	animated,
vilka	who; which; that,which,
tillräckligt	sufficient,
utrustning	equipment,gear,
tillräckliga	insufficient,
svenskarna	the swedes,
yttersta	furthest,
dygn	day,
fiskar	fishes,fish,
uppenbarelser	revelations,
berlinmuren	berlin wall,
motståndarna	opponents,
tankar	tank,thoughts,
sak	substance,
san	san,
sam	co,
generation	generation,
konsekvenser	consequences,
argument	argument,arguments,
församlingar	parishs,assemblies,
say	say,
känslan	the feeling,
burundi	burundi,
allen	allen,
turner	tournament,
västberlin	west berlin,
övriga	other,others,
takt	rate,
styrelsen	the board,board,
zoo	zoo,
massa	mass,
förändringen	the change,
föder	give birth,gives birth,
muslimer	muslims,
finlands	finlands,
sekreterare	secretary,
tränare	coach,
knep	tricks,
religionen	religion,the religion,
religioner	religions,
rådets	council,
kontroversiell	controversial,
driva	run,
förändras	changes,
inledningen	the introduction,
ursprung	origin,
fredspriset	peace price,
rykte	reputation,
kvicksilver	mercury,quicksilver,witty zeal,
katekes	catechism,
rött	cane,red,
olagligt	illegal,
axl	axl,
genomförts	out,
beckham	beckham,
dahléns	dahlén's,
sjöss	sea,
antalet	number,the number,
stärkte	strengthened,increased,
slog	hit,
heinrich	heinrich,
beatles	beatles,
kategorimusik	category music,
återvänder	returns,atervander,
egentliga	real one,actual,
platta	flat,
spetshundar	sets dogs,tip of dogs,
ländernas	countries',countries,
artist	artist,
råd	advice,council,
enighet	unity,
översättningen	translation,the translation,
roger	roger,
ljudet	the sound,noise,
varna	varna,
yta	surface,
monark	monarch,
erbjöds	offered,
dagsläget	current situation,
översättning	translation,
spetsen	edge; top,
brännvin	aquavit,
snabbare	rapid,faster,
behovet	need,the need,
up	i[,
nederbörden	precipitation,the precipitation,
skärgård	archipelago,cutting garden,
talman	speaker,
personlighet	character,
enhetlig	single,
utgörs	is,make up,
förvaltning	administration,
källa	source,
kritiserade	criticised,
begränsningar	limits,
upplever	experiencing,
kontrakt	agreement,contract,
kilometer	kilometers,
revolutionär	revolutionary,revolutions,
amerikanskt	american,
anledningarna	reasons,
screen	screen,
fynd	finding; finds,findings,
antika	ancient,
amerikanske	american,the american,
awards	awards,
inverkan	influence,effect,
amerikanska	u.s.,american,
mariette	mariette,
basisten	bassist,
skönlitteratur	fiction,
nationell	national,
s	s,
rekord	record,
mani	mani,mania,
tillsätts	added,appointed,
långsammare	more slowly,slower,
upproret	revolt,rebellion,
hamnade	ended up,
drogs	was,
därtill	thereto,
farfar	grandfather,
airlines	airlines,
dödsfall	death,deaths,
luft	air,
cupen	cup,
lidit	suffered,
förr	sooner; past,sooner,
formen	the form,
formel	formula,
arabiska	arabic,arabian,
tillåter	allows,allow,
tillåtet	allowed,
pernilla	pernilla,
former	forms,
landskapen	the landscapes,landscapes,
samling	concentration,collection,
representativ	representative,
friska	healthy,fresh,
situation	situation,
föregångaren	predecessor,
peruanska	peruvian,peruan,
förlängning	overtime; extension; prolongation,
startar	start,
bron	bridge,the bridge,
tillåtelse	permission,allowed,
sammanfaller	coinciding,coincides,
beteckna	denote the,denote,
ohälsa	disorders,
världsbanken	world bank,
försäkra	insure,
träffat	met,
ärftliga	genetic,
otto	otto,
träffas	meet,reached,
oceanen	ocean,
ekologi	ecology,
sägas	is said (to be),
lindgrens	lindgren's,lindgrens,
förkortning	abbreviation,
senator	senator,
personlighetsstörning	personality disorder,
måla	grinding,
tillfälle	time,
gestalter	beings,figures,
avser	regards,regard,
ifrågasatt	question,
iraks	iraq,
gudomliga	divine,
förluster	losses,
bokförlaget	publisher,
berättelse	tale,story,'s re,
koncentration	concentration,
spårvagnar	trams,saving carriages,
psykologisk	psychological,
likheter	similarities,similarity,
resa	travel,
libyen	libya,
förlusten	loss,
judarnas	jews,
kastar	castes,throws,to throw,
unika	unique,
helige	holy,
miljon	million,
instrument	intrument,
körberg	körberg,
infördes	introduced,
unikt	unique,
heligt	holy,
störst	most,
snart	soon,
vinkel	angle,
dark	dark,
regim	regimen,regime,
unesco	unesco,
litteraturen	literature,
gotlands	gotland,
skadade	wounded,
stammar	strains,stutters,
vattenånga	steam,
stupade	fallen,killed,
fossila	fossilized,fossil,
intet	nothing,no,
nämnas	mentioned,worth mentioning,
what	what,
ansvar	responsibilities,
ursprungsbefolkning	indigenous,
ekman	ekman,
kännedom	knowledge,
närheten	near,the vicinity,
björn	björn,bear,
föreslog	suggested,
institutionerna	institutions,
ddr	ddr,
exil	exile,
cannabis	cannabis,
atomkärnor	nuclei,nuclear particles,
ingående	input,
västerås	västerås,
katolsk	catholic,
långstrump	hose drumstick,
jacksons	jackson's,
nivån	level,
medlemsstater	member,member states,member-state,
stone	least,
organisationen	the organization,
ace	ace,
väldet	empire,
populationen	population,
befinner	is,placed; situated; positioned; are,
populationer	populations,
organisationer	organizations,organisations,
visst	specific,certain,
billboardlistan	billboard list,bilboardlist,
upplevelser	experiences,
ronden	round,
bryts	breaks,
nationalencyklopedin	national encyclopedia,the national encyclopedia,
image	image,
säkerhetsrådet	security,
partiet	the party,
bryta	break,
partier	parties,
bergen	mountains,
striderna	the battles,fighting,
förintelsen	holocaust,
philadelphia	philadelphia,
evangeliska	evangelical,
söker	searches,seek,
hel	full,(whole) lot (of),
hamnen	harbour,the harbour,
sover	sleep,
hänger	hanger,
hänvisning	reference,
dagen	day,
complete	complete,
bevarat	preserved,
bevaras	are protected,preserved,
mick	mike (microphone),
kontroverser	controversies,
språkliga	linguistic,language compatible,
bevarad	preserved,
rush	rush,
uppträdande	conduct,
jamaicas	jamaicas,jamaica's,
hexadecimalt	hexa-decimal,hex,
utmed	along,
vinkeln	angle,the angle,
afrodite	aphrodite,
förbundsstat	federal,federal state,
regimer	regimes,
krona	crown,
ac	ac,
ad	ad,
tunisien	tunisia,
gustafs	gustafs,
am	am,
bronsåldern	bronze age,the bronze age,
as	as,
beordrade	commanded,
håll	hold,
väsentligt	substantially,
förhistoria	prehistory,
federala	federal,
riktningar	directions,direction (-s),
svårt	black,difficult,
svåra	answering,difficult,
avslöjade	revealed,
såsom	such as,like,
värmlands	varmlands,värmlands,hot countries,
koppar	copper,
gifte	married,
medverkan	participation,
kvarstod	remained,
kategorisvenskspråkiga	category swedish-speaking,
terra	terra,
medverkat	participated,
värd	host,
terry	terry,
vanliga	regular,
forntida	prehistoric,
kommunen	municipality,
kommuner	municipalities,local,counties,
århundradena	centuries,
nelson	nelson,
omgivningen	the surrounding,
original	orignal,
renässans	renaissance,
känslor	music,
släppt	self-indulgent,
släpps	released,(is) released,
elektron	electron,
koloniserades	is colonized,
anpassning	adaption,adjustment,
kammare	chamber,
års	year,years,
 kmh	kmh,
norr	north,
skogarna	forests,
pojkvän	n/a,boyfriend,
ty	for,
tv	tv,
romanen	novel,
nederbörd	precipitation,
to	to,
romaner	novels,
th	th,
nord	north,
te	tea,
ta	to,
ghana	ghana,
telefonen	phone,
strand	beach,
utländsk	foregin,foreign,
ensamma	alone,
djurarter	species,
sauron	sauron,
muslimska	muslim,
utsåg	appointed,
sand	sand,sandy,
siffrorna	figures,the numbers,
smala	narrow,
harry	harry,
sann	true,
språkbruk	parlance,language,
döttrar	daughters,
samoa	samoa,
synd	sin,
dödsstraff	death penalty,
utökade	expanded,increased,
vägnät	network,
skede	stage,
givaren	the giver,dealer,
richard	richard,
delen	part,
soldater	soldiers,
islams	islams,
leif	leif,
gjorts	made,
hänsyn	light,
full	full,
gruppen	the group,group,
själen	the soul,
arkeologiska	archaeological,
november	november,
legend	legend,
äventyr	adventure,adventures,
hindra	prevent,
traditionella	traditional,
känsliga	susceptible,
traditionellt	traditional,
social	social,
action	action,
oftare	more,
varelser	creatures,
juridiska	legal,
vid	in,by,at,
ordinarie	permanent,regular,
vin	wine,
juridiskt	legally,juridical,judicial,
vis	vis,
kuiperbältet	kuiperbaltet,
vit	white,
spelaren	the player,
skapa	creating,
biskopen	bishop,
mors	mother,mothers,
underordnade	subordinate,subordinates,
sitter	serve,
presenterades	presented,
rhen	the rhine,rhine,
dödligt	deadly,
mora	mora,
bevis	certificate,
mord	murder,
ragnar	ragnar,
berättade	told,
uppskattas	is appreciated,estimated,
uppskattar	estimates,
schweiz	switzerland,
undergång	destruction,
socialt	social,
medelklassen	middle class,
science	science,
monoteistiska	monotheistic,
sociala	social,
morgan	morgan,
studenter	students,
läkaren	the doctor,
samväldet	commonwealth,
sikt	run,
nordvästra	northwest,
skadliga	harmful,deleterious,
staten	state,
mellersta	middle,the middle,
states	states,
stater	states,
spansk	spanish,
järnvägsnätet	rail,
vägnätet	road network,
hugo	hugo,
ansetts	considered,
uppnått	met,
lejon	lion,
retorik	rhetoric,
brett	broad,
produktionen	production,the production,
referens	reference,
lanka	(sri) lanka,
köpte	bought,
barnens	children's,the child's,childrens,
komplext	complex,
pucken	the puck,
komplexa	complex,
utvidgning	enlargement; expansion,enlargement,
hållit	held,
nationerna	the nations,nations,
blommor	flowers,
trade	esterified,
östblocket	east block,the eastern bloc,
kvinnors	women,
aktiviteter	activities,activity,
anställda	employed,
vietnamkriget	vietnam war,
känsla	feeling,sense,
alla	all,
högskola	college,
protestanter	protestants,
caesars	caesars,
miljön	environment,
termen	the term,term,
filip	filip,
alls	all,
få	have; make; few,
stadshus	town hall,city hall; town hall,
isaac	isaac,
samhällets	of society,
berömda	famous,forceps,
inleda	initiate,
sträckor	distances,
privilegier	privileges,
produceras	produced,
passagerare	passengers,
grekisk	greek,
introducerade	introduced,
producerade	produced,
olycka	incident,accident,
intåg	entry,advent,
budskap	message,
målning	painting,
graviditet	pregnancy,
blodet	the blood,blood,
denna	that,
härrör	derived,
enstaka	occasional,single,
populärt	popular,popularly,
sydöst	south east,
doser	dose,
populära	popular,
blues	blues,
förespråkade	advocated,
kretsen	the order,circuit,
finner	found,finds,
uppfördes	built,
massiv	massive,
omröstningen	vote,the election,
kopplad	connected,
garvey	garvey,
avgick	retired,
research	research,
norska	norwegian,
uppstått	resulting,arised,
sammanfattning	summary,
kopplat	coupled; connected,coupled,
kopplas	connected,coupled,
highway	highway,
sparken	park,gets fired,
stjärnor	stars,
driver	run,drive,
båda	both,bath,
både	both,
kostade	cost,
ålands	Åland island's,the Åland island's,
kärnkraft	nuclear power,nuclear,
poeten	poet,the poet,
teknologi	technology,
definition	definition,
service	service,
turistmål	tourist attraction,
persons	persons,person's,
naturens	nature's,
omfattar	encompass,include,
skolan	school,
w	w,
nivåer	levels,
uppenbarelse	revelation,
principen	the principal,principle,
bidragit	contributed,
kristna	christian,
foten	foot,
skiftande	shifting,
spekulationer	speculations,
såg	see,saw,
gemensamma	joint,
avel	breeding,breed,
liknas	compared to,likened,
tove	tove,
sår	wound,
missade	failed,
läggas	laid,added,
chefen	commendant; commander,
tappade	lost,
zeppelin	zeppelin,
moder	parent,
bidrog	contribute,
obama	obama,
organiseras	organizes,organized,
organiserat	structured,
niklas	niklas,
freud	freud,
organiserad	organised,
video	video,
ägg	eggs,egg,
äga	be,own,aga,
väljer	elects,
avslutade	ended,
inkluderar	includes,
generationen	generation,the generation,
förstörelse	destruction,
inkluderat	including,
ägt	taken,
ägs	is owned,(is) owned,owned,
astronomin	the astronomy,astronomy,
visats	demonstrated,
framåt	forward,forth,
varianten	version,variant,
norstedts	norstedt's,collins,
kongokinshasa	kong kinshasa,democratic republic of the congo,congo kinshasa,
varianter	variants,varieties,diversities,
arabisk	arabic,
sträcker	stretches,
sydostasien	southeast asia,
brooklyn	brooklyn,
arter	species,
utsattes	subjected,were exposed,
cover	cover,
kanalen	channel,
kanaler	channels,
arten	species,
mesopotamien	mesopotamia,
golf	golf,
omfattade	included,
falska	fold,false,
presidentens	the president's,the presidents,
detalj	detail,
karaktär	character,
falskt	false,
richmond	richmond,
framgångar	successes,success,
existensen	existence,
betydelser	meanings,
jämföra	compare,
befolkningstätheten	population density,n/a,state of the population,
betydelsen	the meaning,
jämfört	compared to last,compared (to),
karakteristiska	characteristic,
gratis	free,
evolutionen	the evolution,
tekniken	techinque,art,
tekniker	technician,
erkännande	recognition,
victoriasjön	victoria lake,lake victoria,
tanken	the thought,
ledare	conductors,
bytet	the exchange,
populärmusik	popular music,pop music,
kill	kill,kill found,
river	tear,
påverkan	influence,
någon	someone,
nietzsches	nietzsche,nietzsche's,
ses	be,are seen,
ser	see,sees,
förhöjd	elevated,
sex	six,
sed	sed,thirst,
psykologiska	psychological,
uppkomsten	onset,
moçambique	mozambique,
järnväg	railroad,rail,
sen	then,
något	any,
nations	nation,nations,
institutet	institute,
församlingen	parish,congregation,
guinea	guinea,
neutralitet	neutrality,neutral,
fission	fission,
kejsarens	emperors,
stärkelse	starch,
alqaida	al-qaida,
rita	paint,draw,drawing,
europe	europe,
europa	europe,
giftermål	marrige,
avvikelser	deviations,
medvetet	conscious,
stadsdel	district,
medborgerliga	civil,
demografiska	demographic,
forskare	researchers,
bästa	the best,best,
förändring	alteration,change,
messias	messiah,
stå	stand,
halmstads	straw city,
kopia	copy,
samma	same,
transeuropeiska	transeuropean,
upprättades	was established,establish,
olle	olle,
kriser	crises,
church	church,
allierade	allies,
decennium	decade,
sommaren	summer,the summer,
pressfrihetsindex	press freedom index,
väntade	expected; were waiting,waited,
tillväxt	growth,
potentiellt	potential,
kyrilliska	cyrillic,
idén	the idea,
starkt	strongly,
pågår	(in) progress,
föranledde	led,
beskrevs	described,
skönhet	beauty,
fire	fire,
mind	mind,
taube	taube,
hovrätten	court of appeals,the court of appeal,
fritz	fritz,
uppleva	experience,
fritt	free,
euron	euro,
systematik	systematic,
handling	action,
framträder	stand out,
projekt	project,
budget	budget,
individerna	the individuals,
brottslighet	criminality,crime,
pressen	press,
arbete	work; labor,
von	von,
teoretisk	theoretical,
erkänna	recognize,
lokaler	facilities,studios,
korruptionsindex	corruption perceptions index,corruption index,
kritiker	critiques,
barney	barney,
gärning	deed,
möjlighet	oppertunity,
barnet	child,
skalet	the shell,
högste	chief,highest,
barnen	children,
arméer	armies,army,
kritiken	criticism,the criticism,the critique,
laddning	charge,
kategoriavlidna	category deceased,
snarare	rather,
republiken	the republic of,
republiker	republics,
skapade	created,
debatten	debate,the debate,
kring	around,
ledarskap	leadership,
fyra	four,
vargar	wolves,
euro	euro,
normala	normal,
phil	phil,
normalt	normally,normal,
person	person,
johan	john,johan,
kontakter	contacts,
finansiellt	financial,
konkret	concrete,
tunnelbana	subway,
släppas	released,be released,
telegram	telegram,
stockholms	stockholm,
finansiella	financial,
kontakten	conntact,the contact,
mandat	mandate,
fascistiska	fascist,fascistic,
lady	lady,
festivalen	festival,the festival,
nordväst	north west,
festivaler	festivals,
jönssonligan	jönssonligan,jonssonligan,
tomas	tomas,
australia	australia,
format	shaped,format,
turnéer	tours,
teologiska	theological,
melker	melker,
avvisar	reject,
skara	city in south-central sweden (uppland),
samarbete	collaboration,co,
ivar	ivar,
västsahara	western sahara,
samarbeta	co,cooperate,
funnit	found,
skarp	crisp,
utlösa	trigger,
informationen	the information,
alexandra	alexandra,
evangelierna	the gospels,
vojvodina	voyvodina,vojvodina,
lenin	lenin,
saknar	lack(-s),
saknas	missing,
användbar	useful,
utvecklades	developed,(was) developed,
avskaffade	abolished,absolished,
nåd	mercy,grace,
läste	read,
öka	oka,increase,increasing,
brasilianska	brasilian,
turnerade	toured,
religion	religion,
riksförbundet	national association,
säger	claims; says,
be	be,
norra	north,northern,
ugandas	of uganda,uganda,
västra	vastra,
bl	short of "bland" - in the context: bl. a (bland annat) = among others,
bo	living,
bk	bk,
engelska	england,
bokstav	letter,
ordning	system,
santa	santa,
by	by,
källor	source,
ideologin	ideology,the ideology,
bosättningar	settlements,
soldaterna	soldiers,
gemenskaperna	communities,community,
aggressiv	aggressive,
stuart	stuart,
fungerande	effective,
papper	paper,
texterna	text,
inte	not,
clinton	clinton,
colorado	colorado,
syret	the oxygen,oxygen,
hemingway	hemingway,
kravet	requirement,
spridas	spread,disseminated,
kraven	the demands,requirements,
popsångare	pop singer,
uppkallad	named,
orsaken	cause,
förlaget	publisher,
konstantin	konstantin,
veckor	weeks,
kategorimusikgrupper	category of music groups,
dröja	wait,
utbröt	broke out,
samerna	sami,the lapp,
knuten	tied to,knot,
fattigdom	poverty,
förbindelse	connections,connection,
européerna	europeans,
poster	positions,post offices,
rörlighet	movement,
pastor	pastor,
begreppen	the terms,
begreppet	the term,term,
posten	post,the position,
atom	atom,
kritisk	critical,
lovade	promised,
lina	lina,
dröm	syndrome,
fader	father,
cia	cia,
ut	out; up,out,
drogmissbruk	drug abuse, substance abuse, drug addiction,
förekom	ods,was,
ur	from,
distrikt	district,
uk	uk,
erics	erics,
översvämningar	flooding,floodings,
nämner	mentions,names,
dog	died,
diverse	some,miscellaneous,
utbyggt	develpoed,built,
makedonska	macedonian,makedonish,
nationalism	nationalism,
inblandning	incorporation,involvement,
matematiken	mathematics,
händelsehorisonten	place else horizon,
läsare	readers,
värld	world,
edwards	edwards,edward's,
são	sao,
skrivits	down,
innehåller	contains,
nordafrika	north africa,
innehållet	content,
matematiker	mathematician,
upplaga	edition,uppalaga,submission,
individuella	individual,
besegra	defeat,
dominerades	was dominated,dominated,
radikala	radical,
djurgårdens	djurgården's,
ägnar	dedicated,
slås	beat,slas,
land	country,
passagerarna	passengers,
sällskap	company,
symtom	symptoms,
härstammar	derived,
texten	text,the text,
sawyer	sawyer,
texter	texts,
inspelning	recording,
persbrandt	persbrandt,
släpptes	released,
alltför	all too,way too,
bakåt	reverse,
dyraste	most expensive,
hamnar	ports,
hamnat	got,ended up,got in to,
listade	listed,
dancehall	dance hall,
sent	late,
garden	garden,
märken	brands,sign,
kedjan	chain,the chain,
palestinier	palestinians,
kommunistiska	communist,
flöde	feed,
drogen	the drug,drug,
känner	knows,know,
överleva	survive,survival,
tillhörande	associated,belonging (to),
tro	believing,
påverka	impact,
harbor	harbor,
eva	eva,
tre	three,
romerska	roman,
romerske	roman,
opinionen	opinion,
leonardo	leonardo,
bolsjevikerna	bolsevikema,bolsheviks,the bolsheviks,
natur	nature,
regelbundna	regular,
ställde	stood up,asked,
årtionden	decades,
hyde	hyde,
legitimitet	legitimacy,
victor	victor,
antog	adopted,
index	index,
expressen	expressen,
anton	anton,
praktiken	effectively,practice,practically,
indiens	indias,
suveräna	supreme,sovereign,
möjliggör	enables,
birk	birk,
indian	indian,
ledande	conductive,leading,
stadskärna	city core, city center,
led	step,
lee	lee,
upphovsrätten	copyright,
sålunda	thus,
leo	leo,
les	les,
lev	lev,
hälsa	health,tell (him i said hi),
talang	talent,
motorvägarna	the highways,
tegel	brick,
titanic	titanic,
anländer	arrive,arrives,
tillkom	hold back,
insulin	insulin,
opinion	opinion,
artisterna	artists,
huvudvärk	headache,
förlora	lose,
oxenstierna	the oxenstierna,oxenstierna,
mening	meaning,sentence,
indianerna	indians,
anatolien	anatolia,
andreas	andreas,
sekulär	secular,
illegal	illicit,
hemlig	secret,
elever	students,
godkänna	approve,
klaviatur	keyboard,
orkester	orchestra,
projektet	project,
herbert	herbert,
existerade	existed,existing,
författning	constitution,
samspel	interaction,
ytterst	highly,
överlevande	survivor; survivors; surviving,over living,
villor	villas,
edwall	edwall,
lokalt	locally,
bidraget	grant,
advokat	bar,lawyer,
ortodoxa	orthodox,
lokala	local,
peka	point,
gustafsson	gustafsson,
upprätthålla	keep up,maintaining,
process	process,
klassisk	classic,
etta	first,
high	high,
tryckta	printed,
hercegovina	herzegovina,
sydöstra	the southeast,
föregående	preceeding; previous,previous,
halmstad	halmstad's,halmstad,
frågor	questions,
saknade	lacked,
frånvaro	absent,
övergrepp	assult (-s),abuse,
latinska	latin,
delas	divided,
delar	proportions,
delat	shared,divided,
sydvästra	southwest,
kriminella	criminal,
gunwer	gunwer,
profeten	the prophet,
insatser	action,
regeringsmakten	govermental power,government power,
platt	flat,plate,
väckt	brought,woken,
slutsatser	conclusions,
gitarr	guitar,guitarr,
element	elements,
lundgren	lundgren,
slutsatsen	concluded,the conclusion,
napoleons	napoleon,napoleon's,
byggnadsverk	building,construction,
borde	should,
handboll	handball,
diskar	disks,
houston	houston,
möjligt	possible,
hårdast	the most,hardest,
universiteten	universities,the universities,
delad	divided,
hunnit	had,had time to,
byttes	was exchanged,
universitetet	university,
stundom	sometimes,
möjliga	possible,
solvinden	the solar wind,solar wind,
västerbottens	västerbottens,västerbotten's,
eliten	the elite,
uppdelat	divided,
tecknet	the sign,
uppdelad	split,
sänts	sants,sent,
beståndsdelar	constituents,
ovanlig	uncommon,
konkurs	bankruptcy,
bekant	known,
bryter	breaks,
dock	nevertheless,however,
utgår	deleted,
rotation	rotation,
huvuddelen	main part,
sönder	probes,
peking	peking,
kapten	captain,
intressen	interests,
fortsätta	remain,continue,
smallwood	small wood,
överföras	transfer,
intresset	interests,the interest,interest,
klar	done,
bay	bay,
etymologi	etymology,
matrix	matrix,
borderline	borderline,
trycktes	printed,
utbildad	educated,
enskilda	individual,
umgänge	company,intercourse,
kapitalismens	capitalism,capitalism's,
marxistiska	marxist,
fram	out,
undertecknades	signed,
redskap	tool,
egenskaperna	the qualities,properties,
mötte	met,
statschef	head of state,
underverk	wonder,
uppe	top,up,(on) top, up, above,
lundin	lundin,
förts	brought,
dubbel	double,
förändra	change; alter; replace,change,
kompositör	composer,
krävt	taken,
våldsam	violent,
krävs	needs,
david	david,
blanda	mix,
profeter	prophets,profets,
helst	rather,
davis	davis,
hussein	hussein,
kräva	require,demand,
skillnad	difference,
åring	year old,
jesus	jesus,
användningsområden	possible use,applications,
schweiziska	swiss,
nordkoreanska	north korean,
studerade	studied,
nationalistiska	nationalist,
system	system,
syster	sister,
hebreiska	hebrew,
tränga	push (aside),cut in,
teatern	theater,
blivit	become,
utbyggnad	addition,
havet	sea,
pristagare	laureate,prizewinner,
konservativ	conservative,
utländska	foreign,
haven	the seas,
visdom	wisdom,
samverkar	co,co-operates,
roberto	roberto,
väsen	being,entity,
reagans	reagan's,
troende	believers,
samverkan	co,
jonatan	jonatan,jonathan,
räcker	enough,
användaren	user,
inre	inner,
förslag	proposal,'proposal,proposed,
kritiskt	critical,
instruktioner	instructions,
mills	mills,
filosofin	philosophy,
sinatra	sinatra,
kritiska	critical,
best	best,
uppträdde	appeared,occurred,
viss	certain,
finsk	finnish,
säkert	securely,
när	when,
nät	web,net(work),
trosbekännelsen	creed,faith of confession,
detta	this,delta,
vardagen	vargaden,
kvinnliga	female,
visa	see,
uppror	rebellion,
jul	christmas,
förutsättningarna	conditions,
medan	while,
framgår	will be seen,is shown,
synliga	visible,
våren	spring,the spring,
bred	broad,
bokstaven	the letter,character,
nordöst	north east,northeast,
synligt	wisible,seen,visible,
uppdelade	divided,
hopp	hopes,
fursten	prince,
östfronten	eastern front,
samisk	samian,sami,
jan	jan,january,
religionens	religion's,
liksom	and,as is,
jah	jah,
jag	i,
skarsgård	cut farm,skarsgård,
ilska	anger,
handla	act; buy; consume,
abba	abba,
parlamentet	parliament,
lägger	lies,add,
fotbollsspelare	football player,footballers,
lucky	lucky,
generalen	the general,
parlamenten	the parliament,
meter	metre,meter,
tidigaste	earliest,
britterna	the brits,
h	h,
pirate	pirate,
iranska	iranian,
rymmer	holds,
guvernör	governor,
myndigheterna	authorities,
debuterade	debuted,
michail	michail,
priser	rates,prizes,
avlidit	perished,
priset	the prize,rate,
kronisk	chronic,
lämplig	suitable,
freddy	freddy,
vietnams	vietnam,
författarskap	the writer,
sjöng	sang,
upprättandet	establishment,
längst	longest,
balansen	balance,the balance,
varning	warning,
kategorisvenskar	category swedes,
finalen	final,
bolivias	bolivia's,bolivia,
strider	strides,conflict,battles,
bilar	cars,
ende	only,
förklaringar	explanations,
kedjor	chains,
islamiska	islamic,
ett	a,one; a; an,
marknaden	market,
beläget	located,base,
fåglar	birds,
norge	norway,
ogillade	disliked,
belägen	located,situated,disposed,
utövade	exerted,exercised,
tätbefolkade	populated,
ekvatorn	equator,
religiösa	religious,
botten	the base,
co	coli,
dör	dies,
ca	cirka,approximately,
mengele	mengele,
cd	cd,
sannolikhet	probability,
död	death,dead,
bröllop	brollop,wedding,
stabila	stable,
musikvideo	music video,
dök	appeared,dove,turned,
antal	number of,
jussi	jussi,
keltiska	celtic,
moraliskt	moral,
överallt	in all,overall; everywhere,
kombination	combination,
växt	plant,
genetik	genetics,
moraliska	moral,
antas	is required,expected (to),
antar	adopting,adopt,
typisk	typical,
frågorna	questions; issues,
molekyler	molecules,
tvungna	forced,forced to,
puerto	puerto,port,
atlanta	atlanta,
mandatperiod	term,term (of office),
långsamma	slow,
erhöll	obtained,acquire,
rikets	its,the kingdom's,
demokrati	democracy,
vd	ceo,
ondskan	evil,
förlopp	process,pattern,developments,
omnämns	mentioned,
vi	we,
kurdistan	kurdistan,
vm	world championship,vm,
lust	loss,
flickor	girls,
föreligger	is,
sitt	its,
slovenska	slovenian,
utfärdade	issued,
tupac	tupac,
armé	poor,
medeltida	middleaged,medieval,
foundationthe	the foundation,
huden	skin,
paulo	paulo,
känd	known,unknown,
terrorism	terrorism,
flesta	most,
ball	ball,
framförde	performed,
anordnas	organised,
anfield	anfield,
sjukhus	hospital,
diabetes	diabetes,
representera	represents,
mänskligt	human,
väger	weight,
vägen	the road,
ledde	resulted,led,
ledda	run (by),
gatan	street,the street,
kontakt	plug,contact,
kiss	kiss,view,
summan	sum,
paul	paul,
pappa	dad,
frånträde	relinquishment,
tolkade	interpreted,
derivata	derivative,
kunder	clients,
nacional	nacional,
frågan	issue,the question,
framtid	future,
förknippad	associated,
motorvägen	highway,
government	government,
ledarna	the leaders,
dess	then,its,
arbetarklassen	working class,
tillverkning	production,
pressas	pressed,
följeslagare	companions,companion,
lät	had,
emma	emaa,emma,
lär	learn,
aktiebolag	limited company; joint-stock company,stock company,
vallhund	herder,
stadsbild	cityscape,
amazonas	amazon,amazonas,
symptomen	symptoms,
högskolan	hogs school,college,
flotta	fleet,
uppskattades	estimated,appreciated,was appreciated,
tackade	said/thanked,
visade	showed,
miniatyr|	miniature,
filmografi	filmography,folmografi,
anarkismen	the anarkism,anarchism,
trotskij	trotskij,trotsky,
lägsta	minimum,
stannar	stop,stays,
transport	carriage,transport,
skriftliga	written,
februari	february,februari,
kolonin	colony,
behandlades	treated,
flitigt	frequent,
tänkandet	thinking,
dags	time,
naturlig	natural,
kollektivtrafik	public transport,
svaga	faint,weak,
fråga	ask,
biologi	biology,
ateism	atheism,
östberlin	east berlin,
svagt	weak,
gandalf	gandalf,
smärta	pain,
vargen	the wolf,
användande	use,use; usage,
kontinenten	the continent,
må	mon,
erövrade	conquered,
blodiga	blooded,
angeles	angeles,
kontinenter	continents,
lysande	brilliant,
solsystemets	solar system,
burma	burma,
anpassade	adjusted,custom,
släpper	release,
upplösningen	dissolution,
sekelskiftet	the turn of the century,
planetens	planet,the planets,
kristus	christ,
mera	more,
varma	hot,warm,
bedöma	judge; decide,assessment,
skola	school,
blå	blue,blah,
fläckar	stain,
bedöms	judged,evaluated,
överbefälhavare	commander-in-chief,supreme commander,
stadium	stage,
radioaktiva	radioactive,
samlingar	collection,
förre	forrester,
indonesien	indonesia,
apollo	apollo,
radioaktivt	radioactive,
svält	starvation,starvations,
återkommer	recurs,will return,returning,
official	official,
volvo	volvo,
stormakt	great power,major power,
monument	monuments,
inrättades	established,were implemented,
distribution	distribution,
ovanför	over,above,
kingston	kingston,
heter	is named,
utnyttjar	using,uses,
utnyttjas	utilized,used,
skilsmässa	divorce,
separerade	separated,
särskild	specific,particular,
banan	banana,
vitryssland	belarus,
sharia	sharia,
brandenburg	brandenburg,
distinkta	distinct,
lutning	closing,angle,
relationen	the relation,ratio,
månaden	the month,
oavgjort	tie,draw,
modernistiska	modernistic,modernist,
bröd	bread,
övergång	transition,
francisco	fransisco,
uttalade	commented; made a comment; spoke about,stated,
fristående	independent,stand-alone,
förhandlingar	negotiations,
syskon	sibling,siblings,
sänker	sinks,
mineraler	minerals,
kommersiell	commercial,
nederländska	dutch,
näsan	the nose,nose,
child	child,
elisabeth	elisabeth,
bosniska	bosnian,
representanthuset	house of representatives,
invadera	invade,
preussen	prussia,
konsekvenserna	impact,
smålands	smaland's,
atlanten	atlantic,the atlantic ocean,
bibel	bible,insulin,bilble,
spel	game,
edward	edward,
nervsystemet	nervous system,
ale	ale,
mördade	murdered,
främsta	request,primary,
främste	chief,premier,
geologi	geology,
jacob	jacob,
innefattar	comprises,includes,
slutliga	evenutal,ultimate,
upphörde	ceased,expired,discontinued,
estland	estland,estonia,
jamaica	jamaica,
starkast	strongest,
ständerna	the cities,
sabbath	sabbath,
horn	horn,
chef	head,
alltsedan	even since,since,
förbättringar	improvements,improvement,
eurovision	eurovision,
bakgrunden	background,
vidsträckta	broad,wide; broad,
kraftfull	powerful,
tolv	twelve,
bidrag	contribution,contributions,
vampyr	vampire,
cyklar	bikes,
bidrar	contributes,
petra	petra,
musikalen	the musical,
räddar	saved,
bortgång	passing,death,
pluto	pluto,
norstedt	norstedt,
same	lapp,
begått	comitted,committed,
interna	internal,
studeras	is studied,
studerat	studied,
interstellära	interstellar,
regerande	ruling,
hänvisade	referenced,referred,refer,
förblir	remain,
stoft	dust,
placerades	placed,
akc	akc,
kongressen	congress,
järnmalm	iron ore,
faktiskt	in fact; actually; indeed,really,actually,
läkemedelsverket	medical products agency,medicines work,food and drug administration,
tillsammans	together,
faktiska	actual,
absolution	absolution,
sarah	sarah,
ätten	the dynasty,dynasty,
negativa	negative,
foster	fetus,
negativt	negative,
supportrar	supporters,
ifall	if,
giovanni	giovanni,
fingrar	finger,
riksväg	national highway,
alces	alces,
lissabonfördraget	lisbon treaty,
kurderna	kurdish,
springer	running,springer,
friheten	liberty,
ik	ik,
era	era,
transparency	transparency,
skiljer	differs,is different; differ,
folkmun	popular lore; popularly,
vackra	beautiful,fine,
felaktiga	false,
ekonomiskt	economically,economical,
in	in the context: recorded = spela (in),in,
indien	india,
felaktigt	incorrect,erronenous,
marco	marco,
enhet	unit,entity,
valborg	valborg,
uppmärksamhet	attention,attantion,
solen	the sun,sol,
firas	celebrated,celebrate,
firar	celebrate,
gillar	enjoy; like,
halland	halland,
beach	beach,
sammansatt	compound,
rädd	scared,afraid,
biografer	movie theaters,cinemas,
kategorieuropas	category europe,
lag	act,
koreakriget	korean war,
visste	did,
biografen	the cinema,movie theater,
law	law,
orden	words,
medlemsstat	member state,
vänsterpartiet	left wing party,
lämningar	remains,
massmedia	media,
livets	life,life's,
offentlig	public,published,
arbetslöshet	unemployment,unemplyment,
sovjet	soviet,
inspelningarna	recordings,
blandning	mix,mixture,
bidra	contribute,
straff	penalty,punishments,
lagets	substrate,the team's,
fragment	fragment,
vanligtvis	generally,
ämne	substance,subject,
fredsbevarande	peace,
bana	course,web,
they	they,
spelningen	the gig,the concert,
bank	bank,
huvudartikel	main article,
l	l,
dåliga	poor,bad,
diskuteras	discussed,is discucssed,
knutpunkt	hub,
tendens	tendency,
dåligt	poor,
område	area,
erbjöd	offered,
germanska	germanic,germanian,
voddler	voddler,
däggdjur	mammalian,
rummet	room,
kejserliga	imperial,
lugna	calm,
daniel	daniel,
därav	thereof,
trafik	traffic,
bruttonationalprodukt	bnp,
veta	out,
värdefulla	valueable,
standard	standard,
förmodligen	presumably,
tillbaka	back,
berör	affecting,affect,
ange	set,name,
sprit	liqeur,
väldiga	vast,
professionell	professional,
höll	held,hold,
personerna	people; persons,the persons,
funktioner	functions,features,
önskar	desiring to,
önskan	desired,
statskupp	coup,
ingmar	ingmar,
synnerligen	remarkably; particularly,particularly,quite,
kantonerna	cantons,
begränsas	begransas,
begränsar	limit,
ingen	no,
sång	song,
förklarade	explained,said,
växthusgaser	greenhouse gas,
inget	not,no,
begränsad	limited,
medborgare	citizens,
antisemitismen	antisemitism,anti-semitism,
äter	eat,eats,
militärt	military,militarily,
albert	albert,
kvarvarande	residual,lasting,
persson	persson,
bojkott	boycott,
kraftverk	plant,
källkod	source,source code,
religionerna	religions,the religions,
symboliserar	symbolized,symbolizes,
binda	tying,bond,
kronan	kronan,swedish krona,
sonen	the son,
scener	scenes,
används	use,used,
scenen	stage,
binds	bound,(is) bound,
iron	iron,
minut	minute,
använde	used,
använda	using,
årens	years,
skolorna	schools,the schools,
fåglarna	the birds,
omvandling	transformation,
framtida	future,
koloniala	colonial,
anledningar	reasons,
kalendern	calender,
stavning	spelling,
magnus	magnus,
höjd	height,
sjukvård	health care,healthcare,
aftonbladet	newsweek,the evening paper,
lades	put,
anatomi	anatomy,
närvaro	attendance,presence,
historisk	historic,historical,
verkar	acting,seems,
maiden	maiden,
utställning	display,exhibition,
skansen	forecastle,
fjädrar	feathers,
flygplatsen	airport,the airport,
eviga	eternal,
ägda	owned,
freja	freja,joe,
ägde	tookplace; occured,
bortom	beyond,
läran	laran,
evigt	forever,eternal,
effekten	effect,
damer	ladies,
lewis	lewis,
hinduiska	hindu,
vanligen	usually,typically,
effekter	effeckter,
rankning	ranking,rating,
sättet	manner,way,the way,
 kilometer	kilometer,
sätter	puts,
näring	nutrition,
estetiska	aesthetic,
bevarats	preserved,
kejsar	emperor,
inställning	attitude,
målvakt	goalkeeper,
variera	vary,
do	do,
imperium	empire,
dj	dj,
di	di,
dc	d.c.,
da	da,
stalins	stalin,
watson	watson,
människorna	men,
orolig	worried,
riktningen	direction,denomination,
du	to,you,
dr	doctor,doktor,
peyton	peyton,
offret	the victim,offering,
runt	around,between,
emo	emo,
konst	art,
offren	victims,
tyngre	heavy,heavier,
fågelarter	bird species,
lasse	lasse,
libanon	lebanon,
veckan	weeks,
vanlig	ordinary,common,
utförd	performed,
utföra	perform,out,
förena	combine,unite,combining,
stewie	stewie,
historiens	historys,history's,
utfört	done,
massiva	solid,massive,
djuret	the animal,animal,
fornnordiska	old nordic,
månarna	moons,
fångenskap	captivity,
piratpartiet	pirate party,
materialet	the material,
smaken	flavor,
osmanska	osmanian,ottoman; osmanli,
komplikationer	complications,
we	we,
självständigheten	independance,independence,
intog	seized,occupied,took,
miljö	environment,
jämförelse	comparative,comparison,
huvudsakligen	generally,primarily,
militären	military,the military,
muhammed	muhammed,
startade	started,
kommer	is,
brad	brad,
gruppens	group (-s),group,
målningen	milling,
kännetecken	sign,
thierry	thierry,
fångar	prisoners,
tusentals	thousands,
genomför	implement,
tony	tony,
japans	japan's,
patienten	patient,
tids	time,
lösning	solution,
framträdande	apperance,appearance,
hitlers	hitlers,
patienter	patients,
nära	close,
attacken	attack,
attacker	attacks,assaults,
fest	festival,fest,
juridik	law,
frekvens	frequency,
bulgariens	bulgaria's,bulgaria,
fromstart	starting from,
vagn	wagon,
johansson	johansson,
påstådda	said,alleged,
kupp	kupp,coup,
nordöstra	northeast,
spanjorerna	spaniards,
gärdestad	garden city,
moldavien	moldova,
deltagarna	the participants,
jordbruk	agricultural,
påverkades	affected,
sagor	fairytales,fairy tales,
patent	patent,
datorer	pc,
bergskedjor	mountain ranges,
självt	itself,
utgivna	published,
bunny	bunny,
andelen	the proportion,
platina	platinum,
hann	did,managed to (in a period of time),
saddam	saddam,
balkan	balkan,
sexualitet	sexuality,
delstater	states,
hand	hand,care,
delstaten	land,
hans	his,
bilen	car,
koncentrerad	concentrated,concentration,
aspekter	aspects,
förlorade	lost,
rörelsen	movement,
kyla	cold,
riksdag	parliament,the parliament,
rör	touch, move(-s),touches,
styrkorna	forces,
mamma	mother,
monaco	monaco,
rörelser	movements,
röd	rod,
thc	thc,
skottland	scotland,
gärningsmannen	the offender,culprit,
newton	newton,
kall	cold,
nästan	almost,
goda	good,
enades	agreed,
kalender	calender,
upptäckte	found,
swahili	swahili,
lindh	lindh,
så	so,
påföljande	following,
wright	wright,
havets	the seas,
kvinnan	female,
plasma	plasma,
född	born,
förbättra	improve,
föda	feed,give birth,
rna	rna,
skadorna	damage,injuries,
arab	arab,
indianer	indians,
föds	born,
everton	everton,
picasso	picasso,
hepatit	heptatitis,
acceptera	acceptable,
årlig	yearly,
indelning	classification,
dahlén	dahlén,
samfund	communities,
gandhi	gandhi,
transkription	transcription,transcript,
avsätta	unseat,
born	born,
presidentvalet	presidential election,
bord	table,
kungar	kings,
humor	humor,humour,
territorierna	territories,
purple	purple,
serbiens	serbias,
siffran	number,
vinterkriget	the winter war,winter war,
stadsdelarna	districts,
vägar	paths,
bevara	preserving,
fängslades	imprisoned; jailed, gaoled; incarcerated,jailed,
slovakien	slovakia,
upplösning	resolution; dissolution,resolution,
banker	banks,
olika	different,variety,
samer	sami,
roms	rome's,roms,romes,
karlsson	karlsson,
epicentrum	epicentre,epicenter,
fängslade	imprisoned,
blivande	future,to be,
way	way,
was	was,
war	war,
etablerat	established,
hypotes	hypothesis,
skiljas	separated,
motorvägar	highways,motor,
inträffat	occurred,
partiledare	party leader,
emil	emil,
reser	travels,rise,rises,
studierna	studies,
långvarig	of long duration,long,
träning	practice,
erövra	conquer,
engagerade	dedicated,engaged,committed,
moore	moore,
utomlands	abroad,
tesla	tesla,
efter	after,
bilderna	the pictures,
moln	cloudy,cloud,
toppen	peak,
cellerna	cells,
arkitekten	architect,the architect,
förmåga	ability,
janukovytj	janukovytj,
möte	meeting,
arkitekter	architects,
götaland	gotaland,
konservatism	conservatism,
femton	fifteen,
tottenham	tottenham,
reglerar	controls,
regleras	controlled,regulated,is regulated,
rätter	dishes,
hemma	home,
omgivande	surrounding,
rätten	right,the court,
solens	solar,
uppfanns	was invented,
tenderar	tend,
datum	date,
förklaringen	the explanation,statement,
lider	suffering,suffers,
utkämpades	fought,
förhistorisk	forhistorisk,prehistorian,
afrikaner	africans,
heller	neither; nor,
rådet	the council,council,
igelkott	hedgehog,
vänder	vander,face,
division	division,
hannah	hannah,
uttrycka	express,
enskild	single,
hannar	males,
vegas	vegas,
uttryckt	expressed,
avbröts	canceled,interrupted,
enskilt	individually,single,
salvador	salvador,
stycken	pieces; parts,pieces,
gud	god,
nedsatt	impaired,reduced,decreased; diminished,
datorspel	video game,computer game,
hisingen	hisingen,
frigörs	released,
säte	sate,
idéer	ideas,
templet	the temple,temple,
revolution	revolution,
cosa	cosa,
engagerad	dedicated,
invandrade	immigrant,
sköttes	handled,
mål	mal,
formellt	formally,
motsatte	opposed,
stimulera	stimulate,stimulating,
motsatta	opposite,
tidig	early,
ingick	were included,was,
uniform	uniform,
fastigheter	properties,
utspelar	set,
versionen	edition,
gener	genes,
muslim	muslim,
lärde	learned,
marxismen	marxism,the marxism,
påstår	states,claims,asserts,
genen	the gene,
oerhört	extremely,
tillträde	access,
antarktiska	antarctic,
flames	flames,
sistnämnda	last,
avsnitten	chapters,
franklin	franklin,
ponny	pony,
history	history,
vinnare	winner,
ekr	ad,
churchill	churchill,
dåtidens	past times,yesterdays,that time,
extra	extra,
vapnet	the weapon,the weapon; escutheon; coat of arms; arms; badge,
spridit	spread,
vapnen	weapons,
förteckning	label,
fbi	fbi,
presenterar	present,
upprättade	established,
äktenskapet	marriage,
territorier	territories,
stabilitet	stability,
live	live,
regel	rule,
territoriet	territory,
omvärlden	world,
överhuvudtaget	in general,
fransmännen	french,
parallellt	at the same time,parallel,
club	club,
rivalitet	rivality,rivalry,
snabbt	fast,
enda	only,single,
parallella	parallel,
zarathustra	zarathustra,
ämnena	subjects,the elements,
närmar	closing,
kolonialismen	colonialism,
kejsardömet	empire,
snabba	rapid,fast,
ibm	ibm,
ibn	ibn,
interaktion	interaction,
frukt	fruits,
can	can,
heart	heart,
nobels	nobel's,
abort	abortion,
uppstår	occur,
genomgått	passed,
judendomen	the judaism,judaism,
pojke	boy,
betydelse	eea,
kopplingar	connections,
alger	algae,
southern	southern,
riktlinjer	guidelines,
framgångarna	the successes,
gräns	limit,border,
ungern	hungary,
förutsättning	provided,
flyttat	moved,
benny	benny,
michel	michel,
ukrainska	ukrainian,
rekordet	record,
maktens	the powers,forces,
ingripa	interfere,act,
ganska	fairly,
respektive	respective,
generalguvernören	governor-general,governor general,
fält	field,
skabb	scab,scabies,
levde	survived,
därifrån	from thence,from there,
yngre	younger,
varav	which,
halt	content,stop; level,
varar	lasts,
chelsea	chelsea,
nog	enough,
författarna	writers,
förvaras	is stored,
komponenter	components,
terrorismen	terrorism,the terrorism,
jorden	the earth,
nou	nou,
rakt	straight,
now	now,
dödsstraffet	capital punishment; death penalty,the death penalty,
uppgörelse	agreement,
frihet	freedom,
språk	language,
främmande	undesirable,foreign,
antyder	indicates,
stockholm	stocholm,
januari	january,
drog	pulled,drug,
aspergers	aspergers,
em	em,european championship,
sektorn	sector,
citat	quote,
eg	ec,
utbrett	widespread,
spåra	track,trace,
strålningen	the radiation,
ex	eg,ex,
kroatiska	croatian,
kant	kant,edge,
effekterna	the effects,effects,
ep	ep,
er	you,your,
teorier	theories,
återkommande	recurring,
stallone	stallone,
hellre	rather,more preferably,
koffein	caffeine,caffein,
genetisk	genetic,
skära	carve,
marino	marino,
betraktades	considered,
sven	sven,
british	british,
domen	judgment,verdict; judgement,
linné	linen,linneus,
allmänheten	public,general public,
arbetsgivare	employers,
skådespelerska	actress,
förändrats	changed,
ring	ring,
xv	xv,
bergqvist	bergqvist,
våglängder	wavelengths,
konungarike	kingdom,
desmond	desmond,
svenske	swedish,
sheen	sheen,
länder	states,countries,
dessutom	moreover,
satsningar	investments,resources,
spelningar	gigs,
nödvändig	essential,
fascisterna	the fascists,the facists,
delats	divided,been awarded,
television	television,
europeisk	european,
sidorna	the pages,pages,
utbyggda	expanded,expand,
ändrades	changed,was,
kloster	monastery,
grundad	founded,based,
statsminister	prime minister,
faktor	factor,
kairo	cairo,
grundat	founded,based,
grundar	bases,
grundas	based,
anger	indicates,
anges	is put at,
befolkningstillväxt	population growth,
hjälp	help,
hör	include,belong,hears,
skär	skerry,
fortsatte	continued,
fortsatta	continued,
etiopiska	ethiopian,etiopian,
bönor	beans,
hög	high,
skäl	reasons,
kategoriorter	category visited,
numera	now,
successivt	progressively,
egentlig	actual; factual; real,
bekostnad	detriment,expense,
dvärgar	dwarves,
glödlampor	lightbulbs,filament,
sagan	story,
lyfter	lift,
norrmän	norwegians,
nordligaste	northermost,
parlamentets	the parliament's,parliament,
runda	round,
orsaka	cause,
skapats	was created,
doktor	phd,doctor,
kyrkorna	churches,
nazisternas	the nazi's,nazi,
marocko	morocco,
teori	theory,
perfekt	perfect,
mannens	man's,
byggda	constructed,
varmblod	warmblood,warm-blooded,
adolf	adolf,
billiga	cheap,
himmel	heaven,
epoken	epoch,the epoch,
dagbok	diary,log,
mörk	dark,
sydligaste	southernmost,
uppståndelse	resurrection,
mörker	darkness,
samuel	samuel,
gudarnas	gods,god's,
ambitioner	ambitions,
folkomröstning	referendum,
marxistisk	marxist,marxistic,
tävla	compete,
handlingar	actions,
gymnasiet	high school,gymnasium,
facupen	fa cup,
tvingade	forced,forcing,
retoriska	rhetorical,
storstäder	cities,
tillfällig	temporarily,
osbourne	osbourne,
övergången	transition,the transition,
katastrofer	disasters,
depressionen	depression,
uppbyggd	structered,
konstaterade	concluded,established,
ladin	ladin,
depressioner	depressions,depression,
israels	israel's,
import	import,
kommunismens	communism,the communisms,the communism's,
katastrofen	disaster,
sträcka	distance,
ronja	ronja,
ordspråk	saying,proverb,proverbs,
männen	the men,men,
utgivningen	release,the release,
verket	board,
verken	plants,
utgavs	published,
comeback	comeback,
samtal	conersation,call,
monicas	monica,monica's,
mona	mona,
bördiga	fertile,
placerad	disposed,
handlar	is,
kristinas	kristina's,crisis thawed,
propaganda	propaganda,
feminismen	feminism,
nils	nils,
comet	comet,
placerar	place,
placeras	placed,
utnyttja	use,
avskaffande	elimination,abolishment,
regeringens	government,
lägenhet	apartment,appartment,
statsreligion	state religion,
riksrådet	riskradet,privy council; council of state; crown council; senate,privy council,
östtyska	east german,
handlande	action,
oliver	olives,
sättas	turn,
sker	is,
oden	oden,
socialdemokrater	social democrats,
dräkt	costume,
observera	note,observe,
utförda	made,
utförde	did,
elvis	elvis,
funnits	found,
konservativa	conservative,
anslöt	joined,
ytan	the area,
uefacupen	the uefa champions league,uefa europa league,uefacupen,
rapporter	reports,
prinsessan	princess,
rapporten	report,the report,
polens	polands,pole,
ordningen	the order,order,procedure,
ändå	spirit,
ansikte	face,
tjeckien	czech republic,the czech republic,
eran	era,
tycker	do,think,
inslag	impact,elements,
finanskrisen	financial crisis,
tänkande	thinking,
behandlade	treated,
kvarter	block,neighborhoods,
kenya	kenya,
västerländska	western,
katalanska	catalan,
helium	helium,
grundade	based,
slaget	type,
långt	far,long,
orsakade	caused,
programvara	software,
media	media,
långa	langa,long,
talmannen	president,speaker of the riksdag,
kromosom	chromosome,
lite	a little,
figurer	figures,
speciella	special,
offensiven	the offensive,
begär	requests,request,
skivbolaget	record label,the record company,
acdc	ac/dc,
målningar	paintings,
omfattas	subject,
speciellt	particularly,
omgående	immediately,immediate,
ekonomisk	economic,
fredspris	peace prize,
skånes	scania's,
erkänd	acknowledged,
erkänt	recognized,
flaggor	flags,
mynning	muzzle,
forskarna	scientists,
skandinaviska	scandinavian,
tydlig	clear,
framgången	success,the success,
samiska	sami,
eleverna	the pupils,the students,
lagerkvist	lagerkvist,
spänningar	tensions,
föreningar	associations,organizations,compounds,
malcolm	malcolm,
lade	laid,seized,
ditt	your,
strävar	striving; aiming (to; for),
irland	ireland,
hovet	court,
stund	while,momentum,
östergötland	Östergötland,
selma	selma,
amy	amy,
fullt	full; fully; completely,
rebecca	rebecca,
symbolisk	nominal,symbolic,
strävan	endeavor,
nationella	national,
skilda	separate,
miniatyr|en	thumbnail,a minature,
skilde	divided,varied,
nationellt	nationally,
t	e.g.,
låga	low,
lågt	low,
präglades	was marked,
stånd	in the context: (make) the war happen,
slår	states,
användbara	useful,
sålts	sold,
indikerar	indicates,
frigörelse	liberation,
bestämd	fixed,
strindberg	strindberg,
utskott	committee,organ,
strålning	radiation,
bestämt	decided,
nsdap	nsdap,
inuti	inside,
växa	growth,grow,
francis	francis,
övertygad	confident,
ideologi	ideology,
jamaicanska	jamaican,
central	central,center,
nordliga	northern,
socialistiska	socialistic,socialist,
torget	square,torget,
bidragen	the contributions,contributions,
efterkrigstiden	the post-war period,post-war,
välfärd	welfare,
klassiker	classics,classic,
transporter	transports,
karriär	career,
area	area,
satsade	invested,bet,
specifikt	specifically,
stark	strong,
start	start,
anställd	employed,
specifika	specific,
likväl	as well,
gånger	times,
hawking	hawking,
sämsta	worst,
gången	time,
traditionerna	traditions,
expeditionen	expedition,
spänner	span,
minne	memory,
engelskan	the english,english,
tidningarna	papers,
minns	remembers,
miguel	miguel,
bilmärke	car make,make of car,
expeditioner	expeditions,
kostar	costs,
kungen	the king,
grammis	grammy,
sveriges	sweden,
godkände	approved,
evenemang	event,
nere	low,
mongoliet	mongolia,
efteråt	afterwards,
trettio	thirty,
you	you,
köper	making,
knä	knees,knee,
expandera	expand,
drift	operation,
bidragande	contributors,
översätts	translate,is translated,
massachusetts	massachusetts,
bandmedlemmarna	band members,
skuggan	the shadow,
tjänare	servant,
handelsmän	merchants,
morgonen	the morning,
färdas	travels,
export	export,
olympiastadion	olympa stadium,olympic stadium,
energikälla	energy source,
öknen	the desert,desert,
loppet	bore,the race,
råvaror	raw materials,wood,
lämpliga	suitable,
påbörjades	commenced; begun,was started,
lämpligt	suitable,fitness,
fästning	fortress,
klorofyll	chlorophyll,cholophyll,
jensen	jensen,
får	can,
verk	work,works,
osv	etc.,
spår	track,
heaven	heaven,
sverige	sweden,
behöver	need,
louis	louis,
mild	soft,
industrialiseringen	indutrialization,industrialization,
koranen	the koran,
rasism	racism,
magdalena	magdalena,
skiva	disc,
fåglarnas	birds,
egendom	property,
kritiserats	critized,
orgasm	orgasm,
markerade	selected,marked,
trupper	troops,
höja	increase,hoja,
tvskådespelare	tv actor,
besöker	visits,
bedrev	conducted,managed,
fjärde	fourth,
förbjuden	smoking,
bernhard	bernhard,
förbjuder	prohibiting,forbids,
sattes	was added,
inblandad	mixed,
förbjudet	prohibited,
irak	iraq,
avbryta	cancel,
genomförde	carried out,
ersättare	alternate,replacement,
observeras	observed,is noticed,is observed,
uttalat	outspoken,
lämna	leave,
uttalas	pronounced,be pronounced,
medarbetare	employees,coworker,
signifikant	significant,
vår	spring,
dyker	dives,
stulna	stolen,
minst	at least,
boxning	boxing,boxing; pugilism,
våg	vague,wave,
kriget	the war,war,
hoppades	hoped,
perspektiv	perspective,
medicin	medicine,
globen	lobe,
nazityskland	nazi germany,
gick	passed,
grunda	found,base,
dalarna	valleys,dalarna,
kritiserat	criticized,criticised,
nukleotider	nucleotides,
avsedd	adapted,intended,
nathan	nathan,
simba	pool,
taket	ceiling,
tillät	distillate,allowed,
etablerad	established,
förlängningen	elongation,forlajgningen,
planen	the field,
trummisen	drummer,
oecd	oecd,
representerar	represents,
teatrar	theaters,
massan	mass,
ryssland	russia,
avled	died,
okänt	unknown,
utökat	expanded,
ständiga	permanent,
latinamerikanska	latin-american,latin american,
inspelad	recorded,
räknar	counts,
räknas	counted,
lagstiftande	legislating,legislation,
ständigt	always,
mördad	murdered,
företeelser	phenomena,
livslängd	life,
fronten	the front,
rapporterade	reported,
paus	pause,paus,
feministiska	feminist,
vistelse	stay,
herrens	lord,
species	species,
zanzibar	zanzibar,
gälla	valid,be valid,
ledger	ledger,
linköping	linköping,
begränsa	limit,
reidars	reidars,
ytterligare	further,additional,
samarbetet	cooperation,the collaboration,
turkarna	turks,
torde	could,should,
fastän	although,
försök	experiments,expirements,
fc	fc,
fd	former,
ff	ff,
samarbeten	collaborations,
stabil	stable,
vattenkraft	water power,hydroelectric power,hydro,
kostnaden	cost,
byggandet	the building,
skivan	disc,
enzymer	enzymes,
allmänna	general,
korset	cross,
kognitiv	cognitive,
segrar	wins,victories,
sänder	transmits,
dream	dream,
nämnts	mentioned,
tillgångar	assets,
helt	completely,
bloggar	blogs,
helgdagar	holidays,
tornen	towers,
hela	full,
kombinerade	combined,
eros	eros,
hundratusentals	hundreds of thousands,
romance	romance,
kompositörer	composers,compositors,
antagits	adoption,
systems	system,
österrikes	austrias,
mahatma	mahatma,
musikalisk	musical,
bytte	changed,changed it's,swapped,
arsenal	arsenal,
konstitutionella	constitutional,
greps	arrested,(was) arrested,
dyrt	a high price,expensive,dearly,
petter	petter,
närmare	further,close to,
märta	märta,
fulla	full,
skrivit	written,wrote,
die	die,
ifk	ifk,
etnisk	ethnic,
neil	neil,
positionen	position,
märktes	labeled,
positioner	positions,
rättvisa	justice,
aktörer	actors,
bodde	lived,
goebbels	goebbels,geobbels,
lungorna	the lungs,
stödet	support,the support,
stöder	supporting,supports,
känna	known,
efternamn	lastname,
utredningen	investigation,the investigation,
heroin	heroin,
delningen	division,
vasas	vasas,
svarade	accounted (for); answered,said,
etnicitet	ethnicity,
skogen	woods,forest,
skilja	differ; differentiate,
förbättrade	improved,
underhåll	support,entertainment,
kung	king,
skiljs	separated,separate,
sändes	was sent,sent,
utvecklats	developed,
synen	the view,sight,
etiska	codes,
elden	the fire,
riksföreståndare	regent,
minoritetsspråk	minority language,
fabriker	plants,factories,
kallat	called,
taggar	spikes,
synes	seems to,apparently,
miss	miss,
rygg	dorsal,
kanada	canada,
kongresspartiet	congress party,
station	station,
parlamentsvalet	election to parliament,parliamentary elections,
nigeria	nigeria,
brittiska	british,
luminositet	luminosity,
läsa	read,
åkte	went,relegated,
lupus	lupus,
förnuftet	the common sense,
tvungen	had,forced (to),
bildande	forming,founding,formation,
växterna	plants,
stora	large,
långsamt	slowly,
einsteins	once a,einsteins,
andersson	andersson,
värden	values,
haddock	haddock,
stiftelsen	foundation,
gren	crotch,
charlotte	charlotte,
bestämdes	was decided,decided,
medeltemperaturen	median temperature,the average temperature,
tvärtom	on the contrary,
nominerad	nominate,nominated,
demokratin	democracy,
vädret	weather,the weather,
grundarna	founders,
henne	she,
liv	life,
herre	lord,master; lord,
avseenden	respects,regard,
mexiko	mexico,
logotyp	logo,logotype,
sektor	sector,
säsongens	season,the seasons,
kan	can be,
bistånd	aid,assistance,
kap	chapter,
fågel	bird,
utgör	constitutes,
kokain	cocaine,cocain,
polacker	polish,
klädd	coated,
räknade	calculated,counted,
recensioner	reviews,
rådde	was,
osäkra	insecure,
ingenting	nothing,
jupiters	jupiter's,jupiter,
möjligen	possibly,
hänvisar	reference,
muslimsk	muslim; muslem,muslim,
svenskans	the swedish language,swedish language,
sanna	true,
justice	justice,
humanistiska	humane,humanistic,
åländska	Åland swedish,aland,
ikon	icon,
lennon	lennon,
darwin	darwin,
ingå	be a part,include,be included in,
dominans	dominance,
arabvärlden	the arab world,arab world,
tillhört	belonged,
gått	gone,passed,
alexander	alexander,
restauranger	restaurants,
avsaknaden	absence,
stadsparken	city park,city ​​park,
vilket	which,
målare	grinders,
x	x,
tolkiens	tolkien,tolkien's,
grunden	base,
allmänt	commonly,generally; public,
maurice	maurice,
tidigare	earlier,before,
ändamål	object,purpose,
grunder	bases,
mörkare	darker,
flyter	float,
direktör	director,
värdet	the value,
pictures	pictures,
lösa	solve,
pjäser	checkers,plays,
löst	dissolved,1st sentence: loosely; 2nd & 3rd: solved,
läns	county,county's,
chansen	chances,
allvar	earnest,serious,
gudomlig	divine,
köket	cuisine,the kitchen,
revolutionen	the revolution,
produkter	products,
lejonet	havskattfskar,
anor	ancestry,lineage; ancestry,
viljan	will,
kyrkliga	religious,from the church,
bott	lived,lived in,
jeff	jeff,
betydde	ment,meant,
scientologikyrkan	the church of scientology,
linux	linux,
sokrates	socrates,
händerna	the hands,
merparten	most,
minskade	minimum period,decreased,
galilei	galilei,
konsensus	consensus,
gestalt	character,figure,
walter	walter,
isolerade	isolated,
budgeten	budget,the budget,
anthony	anthony,
livet	life,
delades	shared,divided,
genomförs	implemented, carried through,conducted,
socialism	socialism,
belgrad	belgrade,
hegel	hegel,
läses	read,is read,
läser	are reading,
diktator	dictator,siktador,
mängden	the amount,
tillfället	time,
slutar	ends,
slutat	left,
kategorikvinnor	category women,
nationalitet	nationality,
klippiga	rocky,
sorter	varieties,types,
bärande	leading,
lagar	laws,
tillfällen	oppertunities,jobs,
kombineras	combined,
staffan	staffan,
kombinerat	combined,
grant	word,
borgerliga	conservative,
deltagande	participation,
sammanlagt	total,
nöd	distress,emergency,
karl	karl,
kombinerad	combined,
grand	grand,
luxemburg	luxembourg,luxemburg,
folkslag	peoples,
bon	bon,
anklagats	accused,
 km	km,
kommunicera	communicating,
förlag	forlag,
seglade	sailed,
armenien	armenian,
svealand	svealand,
fatta	make,to make,
kurdisk	kurdish,
cruz	cruz,
präglad	marked,characterized,
innersta	innermost,
feminister	feminists,
hotell	hotel,
njurarna	kidney,
tortyr	torture,
skal	shell,skin,
inlett	started,ushered in,initiated,
uppfinnare	inventor,
kallblod	draught horse,
taiwan	taiwan,
gänget	the group,gang,
välkända	known,
varuhus	warehouse,
egenskap	ability,seeks,
djur	animals,animal,
bestå	comprise,
återställa	resett,
lika	similar,alike,equal,
gör	makes,
kulturen	culture,the culture,
enklare	easier,simpler,
baserade	based,
unga	young,
läs	read,
immigranter	immigrants,
innan	before,
känslig	susceptible,
releasedatum	release date,
dylikt	such,
koden	the code,code,
criss	criss,
gandhis	gandhi,
terminologi	terminology,
judar	jews,
begärde	called,
mycket	very,much,
kommenterade	comment,commented,
byggnader	structures,
biträdande	assistant,assisting,deputy,
pierre	pierre,
våldet	the violence,violence,
economic	economic,
byggnaden	building,
syndrom	syndrome,
sammanhängande	connective,
världsarvslista	world heritage list,
vilda	wild,
skapar	creates,
slash	slash,
bägge	both,ram,
sarajevo	sarajevo,
run	run,
steg	step,
rum	(took) place,room,
mellankrigstiden	interwar period,
stjärnans	star's,the star's,
offside	offside,
skrivet	written,
benfica	benfica,
freddie	freddie,
führer	fuhrer,
myndighet	authority,
övergick	transended,
linjen	the line,line,
etablerade	established,
fysiologiska	physiological,
refererar	refer (to),reference,
linjer	lines,
edvard	edward,
länderna	the countries,
block	block,
ida	ida,
fåtal	few,
positiva	positive,
ön	the island,
semifinalen	semifinal,
institut	institute,
sprida	spread,
överst	top,at the top; uppermost,
föreningen	association,
fokuserade	concentrated,focused,
ligga	lie,be,
spänningen	voltage,
visat	found,
heritage	heritage,
spridd	wide spread,
ledamot	member,representative,
japanerna	the japanese,
spektrumet	spectrum,
larry	larry,
strukturer	structures,
drabbats	affected,afflicted,
skull	sake,
ute	out,
nyval	new election,
skuld	debt,guilt,
malin	maleic,
trafikerade	frequent,trafficked,
  km²	square kilometre,km2,
politik	politics,policies,
fiske	fishing,
ligacupen	league cup,
tryck	pressure,
ihåg	remember,
metall	metal,
sydkorea	south koreans,south korea,
hårdrock	hard rock,hardrock,
igenom	through,
krigets	war,
sjunde	seventh,
musikens	music,
kategori	category,
relationerna	the relationships,relations,
berättas	(as) told,is told,
rester	residue,residues,
dras	draw,preferred,make (assumptions, references),
drar	drag,
framstående	prominent,
drag	move,
mästare	champion,
kort	short,
resten	the rest,rest,
vindar	winds,
kors	cross,
tillfälligt	temporarly,temporary,
enade	united,
medför	entails,result,
officerare	officers,
tunga	heavy,tongue,
heath	heath,
tillfälliga	temporary,
folkliga	popular,
tungt	heavy,
svt	svt,
dvs	(det vill säga) namely that,d.v.s.,i.e.,
skyskrapor	high rise buildings; sky scrapers,
bonniers	bonniers,
höst	autumn,fall,
placera	position,place,
indiska	indian,
katt	cat,
företeelse	experience; phenomenon; feature,feature,
ge	give,
tänker	thinking,
go	go,
gm	by,
träd	into,tree,
kate	kate,
världsrekord	world record,
baron	baron,
tillhör	belonging to,
toppar	(that) peaks,
dröjde	not until,
sålt	sold,
wave	wave,
rinner	flow,flows,
kommunismen	communism,
försvarsminister	minister of defence,
michael	michael,
utbredning	distribution,
tidszoner	time zones,
jönköping	jönköping,jonkoping,
stift	pin,
akut	acute,urgent,
oklart	clear,
socialdemokratiska	social democratic,
zh	zh,
derivator	derivative,
mussolinis	mussolini's,
honan	the female,
geologiska	geological,
visserligen	although,
söka	search,searching,
börjar	starts to,
börjat	begun to,begun,
svagare	weaker,
kinas	kinase,chinas,
erövringar	conquests,
hansson	hansson,
bjöd	offered,invited,
polen	pole,
gradvis	gradually,progressively,
genombrott	breakthrough,
experiment	experiment,
avancerade	advanced,
valen	the elections,elections,
gasen	gas,
utrikespolitiken	foreign policy,the foreign policy,
bindande	binding,
innerstaden	inner city,
orsaker	causes,
gåva	gift,
eminem	eminem,
uppgick	total,
ryska	russian,
händelser	handelsar,events,
innebandy	floorball,
integritet	integrity,
västerut	west,westward; west,
chans	chances,
överlevnad	survival,
dopamin	dopamine,
uppfinningar	inventions,
avsedda	aimed,intended,
färöarna	the faroe islands,
vuxen	adult,
italienska	italian,
genetiska	genetic,
personen	person,the person,
utdöda	extinct,
coldplay	coldplay,
kunde	could,
stärka	enhance,strengthen; bolster,
jonathan	jonathan,
sjunger	sings,singing,
mexikanska	mexican,
invigningen	inauguration,
huxley	huxley,
misslyckades	failed,
turkiets	turkey's,
debutalbum	debut album,
blod	blood,
släppts	released,
kenny	kenny,
utomstående	outsider,
linköpings	linkopingas,linköpings,linköping's,
beslöt	resolved,decided,
studioalbum	studio album,
talat	spoken,
fördelningen	distribution,
talas	spoken,is spoken,
talar	speaks,speak,
romantikens	romanticism,
tågen	train,the trains,
sovjetunionen	the soviet union,
fälttåg	crusade,campaign,
folkmängd	population,
kronprinsen	crown prince,
oroligheter	unrest,
fara	danger,
uttalet	pronunciation,
svenskar	swedes,
dödlig	lethal,
fart	off,
fars	father's,
utfördes	carried out,was carried out,
ringde	called,
österrikiska	austrian,
säljer	sells,
reagerar	reacts,
absint	absinthe,
encyclopedia	encyclopedia,
kungliga	royal,
kapital	capital,
högtider	feasts,
fungerade	working,
presidenter	presidents,president,
offentliga	public,
förstördes	was destroyed,
någonting	nothing,anything,
offentligt	public,
öarna	islands,
verklighet	reality,
belopp	amounts,amount,sum,
monarken	monarch,
kyrkor	churche,
allting	everything,
filosofiska	philosophical,
konserten	concert,
zagreb	capital of croatia,zagreb,
ägna	baiting,
läror	teachings,
front	front,
konserter	conserts,
dikt	poem,
intäkterna	the revenues,the revenue,
miniatyr|px|den	miniature,
hunden	the dog,dog,
kläder	clothes,
university	university,
räckte	handed,
förmågor	abilites,capacities,
modo	modo,
täcker	attacks,covers,
vilken	what,which,
föreslogs	was suggested,
skog	forest,
globe	globe,
 procent	percent,
stiger	rises,rising,
osmanerna	ottomans,
apartheid	apartheid,
skov	forestry,episode,
skor	shoes,
illa	bad,
flyr	flees,escapes,
entertainment	entertainment,
förutom	except,
upphör	end,
deltagit	participated,
samarbetat	collaborated,
max	max,
solsystem	solar system,
vinter	winter,
torres	torres,
kropp	body,
bilder	pictures,
lycka	happiness,good luck,
bilden	the image,
förstod	understood,
förbund	union,
kommunala	local,
livsmedel	food,
åter	again,
benämnas	named,entitle,entitled,
svart	black,
strida	fight,
tigrar	tigers,
austin	austin,
partierna	portions,
riksdagsvalet	election to parliament,
evans	mr. evans,evans,
minoritet	minority,
önskemål	desire,
peters	peters,
kategorihedersdoktorer	category of honorary degrees,
spaniens	spain's,
attack	attack,
boken	paper,the book,
mao	mao,
dygnet	day,
infaller	falls,
final	finite, final,
nilsson	nilsson,
belgiska	belgian,
hasch	hashish,
emellertid	however,
styrelseskick	form of government,
lista	list,
definierat	defined,
ben	bone,
definieras	defines,
definierar	defining,defines,
arbetade	worked,
inbördes	intermutual,
israelisk	israeli,
ber	ask,asks,
bet	bit,
julian	julian,
kvinnans	female,
hjärna	brain,
bordet	the table,desktop,
varade	duration,lasted,
förra	last,
benämning	name,
visor	songs,
förlorades	lost,
släkt	family,
attackerna	the attacks,
runorna	the runes,
röst	voice,
förblev	remained,
jorge	jorge,
regn	rain,
montana	montana,
kvarstår	remains,
regi	direction,
tyskar	germans,
sändas	broadcast,sent,
överföring	transfer,
skogar	forests,
långtgående	far-reaching,
platon	platonic,
parker	parks,
minska	reducing,
tolkien	tolkien,
fynden	finds; findings,
allvarliga	serious,
försvara	defend,defending,
skedde	was,
passa	fit,
parken	the park,
hade	had,
basen	the base,
baser	bases,
gemensam	joint,common,
härskare	ruler,
förbli	remain,
varit	has been,been,
överlever	survives,
psykologin	psychology,
boris	boris,
klassiska	classic,
inbördeskrig	civil war,
förbjöd	forbade,forbid,
inflytelserika	influential,
klassiskt	classical,classic,
häst	haste,
kämpade	decreased,fought,
karriären	career,the career,
älskade	loved,loved; beloved,
gray	gray,
evolution	evolution,
processer	processes,
tillgång	access,
mohammed	mohammed,
grav	tomb,grave,
gran	spruce,
influensa	flue,
också	also,
kvadratkilometer	square kilometers,
processen	process,the process,
vänt	turned,
produkten	the result,product,
västindien	west india,
förband	units; formations; bound (themselves),bond,
neutralt	neutral,
korea	korea,
stats	state,
tenn	tin,
gotiska	gothic,
staty	statue,
state	state,
företagets	the corporation's,
ken	ken,bank,
högra	right,
ersätta	replacing,
sovjetiska	soviet,
satsa	bet,
benämningen	the name,the designation,
merry	merry,
jobba	work,
utformning	layout,shape,formation,
problem	problem,
tjänster	services,
synvinkel	angle,perspective,
vulkaner	volcanos,
framgångsrika	successful,successes,succesful,
trädde	come into effect,
varierade	varied,
älskar	loves,
utsträckning	extent,
framgångsrikt	successfully,
partiklar	particles,
uppsättning	equipment,
fördelar	share,
fördelas	distribute,distributed,
kategoribrittiska	category: british,
knst	knst,
johans	johan's,johan,
johann	john,
kings	kings,king's,
sammanhang	connection,context,
christer	christer,
liberala	liberal,
sara	sara,
fokusera	focus,
äldre	old,older,
poet	poet,
påminde	reminded,
poes	poe,poes,
pontus	pontus,
vinci	vinci,
övertalade	over spoke,persuaded,
affärer	business,
spanska	spanish,
spaniel	spaniel,
spanien	spain,
humör	temper,
strömningar	tendencies,
kanarieöarna	canary islands,the canary islands,
 meter	metre,
könsorganen	the reproductive organs,
utgjorde	comprised; consisted of,
platons	platon's,plato,platos,
reaktion	reaction reaction,
nordens	the scandinavian countries',scandinavia,nordic,
rysslands	russia's,
feber	fever,
demo	demo,removed,
rättigheter	rights,
nordirland	north ireland,northern,
måleri	painting,
kategorikrigsåret	category war years,
alfabetisk	alphabetical,
revir	turf,territory,
reformationen	reformation tone,
parti	party,
instabil	unstable,
campus	campus,
varmed	whereby,
begav	went,
dickens	dickens,
korrekta	correct,
flygbolag	airline,carriers,
nationens	the nation's,
rankas	ranks,
broder	brother,
införa	introducing,introduce,
eklund	eklund,
nämligen	namely,
spred	spread,
alperna	alps,the alps,
lagring	storage,
flickan	girl,
strömmen	the stream,
i	in,
kärleken	love,
theodor	theodor,
agnostiker	agnostic,agnostics,
onda	evil,
störta	rush,crash,interfere,
sänds	sends,sands,
omkom	perished,
sofie	sofie,
förekommer	occurs,preferred is,
sända	transmitting,send,
sände	sent,
vida	broad,
uppfylla	fulfill,
reducera	reduce,
natt	night,
nato	nato,
kalle	kalle,
titta	see,watch,
jesper	jesper,
katolska	catholic,
utan	without,
sanning	true,truth,
vanligare	more common,
historia	history,
definitivt	unavoidable,definitely,
klassificering	classification,
lincoln	lincoln,
norges	norway's,
fernando	fernando,
page	page,
regeringar	governments,
lager	layer,
kolonierna	colonies,
laget	stroke,
pojkarna	boys,the boys,
library	library,
förlusterna	the losses,loss,
vardagligt	everyday,
förenklat	simplified,
omöjligt	impossible,
skorpan	crust,
peter	peter,
lagen	the law,
moskva	moscow,
skrifter	writings,
kaspiska	caspian,
hyser	has,accomodates,holds,
folkets	folkers,
slott	castle,
alliansen	the alliance,
fanns	was,
förde	led,out,
skriften	no.,
villkoren	the terms,conditions,
hinder	obstacle,barrier,
meddelade	announced,
journal	joumal,jurnal,
reza	reza,
kromosomer	chromosomes,
halvön	peninsula,the peninsula,
småland	småland,
usas	usa:s,u.s.,
keramik	ceramics,
freedom	freedom,
beslutade	resolved,decided,
samlats	solid,
skrev	said,
polisens	police,the police's,
troligen	probably,likely,
synsätt	viewpoint,
hävdade	argued,claimed,
mytologi	mythology,
betydelsefulla	significant,
glenn	glenn,
washington	washington,
räddade	saved,
tendenser	tendencies,
längsta	maximum,
hammarby	hammarby,
djävulen	the devil,
realiteten	de facto,
afrika	africa,
oändligt	infinitely,
distinkt	distinct,distinctive,
cricket	cricket,
north	north,
delstaterna	states,
neutral	neutral,
ho	ho,
hc	h.c.,h.c,
ha	be,have,
he	he,
svarta	black,
fysik	physics,
allierad	allied,ally,
dator	computer,
pippin	pippin,
komiker	comic,comedian,
förslaget	proposition,research team,
hästar	horses,
invandring	immigration,
bitar	bit,pieces,
beatrice	beatrice,
ordbok	glossary,
ibland	sometimes,
erik	erik,
bosättare	settlers,
motsvarar	comparable,corresponds,
diego	diego,
omväxlande	varied,
sänktes	reduced,
moderaterna	the moderates,moderates,
speciell	specific,
jordbävning	earthquake,
hotade	threatened,
vulkaniska	volcanic,
canada	canada,
stat	state,
hittade	found,
revolutionära	revolutionary,
musikvideor	music videos,
stad	city,
musikvideon	music video,
resulterade	resulted,
stan	town,
bly	lead,
hjärnan	brain,the brain,
stam	strain,tribe,
etiken	ethics,
förekomma	be found,
inser	recognize,realizes,
alkohol	alcohol,
blogg	blog,
felaktig	false,error,
andra	other,
fredrik	fredrik,
flest	most,the most,
buddy	buddy,
likaså	also,as well,
upplagan	edition,
kommersiellt	commercial,
kulturell	cultural,
bli	be,
kommersiella	commercial,
gjordes	was,
kristendom	christianity,
östersjön	balticsea,
vasa	vasa,
åstadkomma	provide,
upplysningen	the enlightenment,enlightenment,
kända	known,
kände	felt,
examen	exam,degree,
disneys	disneys,disney's,
försöka	attempt,
chokladen	the chocolate,chocolate,
avståndet	distance,the distance,
sydväst	southwest,
slogs	fought,was,
sexton	sixteen,
dagens	current,
upp	up,
rollfigurer	role figure,
berlins	berlin's,
gator	streets,
neo	neo,
nej	no,
kommissionen	commission,
unescos	unesco,
tänkte	thought,was going to,
new	new,
tätort	conurbation,
ner	bottom,
ort	neighborhood,
med	with,
genomföra	out,
men	but,
drev	pursued,led,
vinden	the wind,
pedro	pedro,
mer	more,
luther	luther,
geografiskt	geographic,
därpå	thereon,
tillverka	producing,
åka	go,
fyllde	completed,filled,
ajax	ajax,
sju	seven,
pilatus	pilate,
geografiska	geographical,spatial,
dra	pulling,pull; (with)draw,
snabbast	fastest,
magnusson	magnusson,
reste	stood,moved,
£m	million pounds,
efterföljare	following,follower,successors,
rosenberg	rosenberg,
reagan	reagan,
inleddes	started,initiated,
fördelning	distribution,
gävle	gävle,
lennart	lennart,
provisoriska	provisional,
rockband	rock band,
oscar	oscar,
ljus	light,
berlin	berlin,
ljud	sounds,noise,
köln	cologne,köln,
flora	flora,
trots	although,
procent	per,
kapitalistiska	capitalistic,
sundsvall	sundsvall,
kanadas	canada's,
erövringen	conquest,
tidskriften	magazine,
abstrakta	abstract,
förväntade	expected,
talets	century,
klitoris	clitoris,
tusen	thousands,
tidskrifter	magazines,periodicals,
vänster	left,
satt	sat,
nobelstiftelsen	nobel foundation,
bonaparte	bonaparte,
avrättningen	execution,
trött	tired,
begrepp	term,
polis	police,
stilla	still,
densitet	density,
orsakas	causes,caused by,
orsakat	caused,
utomeuropeiska	overseas,non-european,
gård	house,
könsorgan	was organ,sex organ,
klarar	handle,
president	president,
orsakad	induced,
indelat	divided,
medföra	bring,result,
indelas	divided,categorized,
indelad	divided,
medfört	led to,resulted,
indisk	indian,
ändra	change,
färdig	pre,
förfäder	ancestors,
fifa	fifa,
centrala	central,
panthera	panthera,
ibrahimović	ibrahimovic,
munnen	the mouth,mouth,
murray	murray,
föreställningar	performances,
helena	helena,
buddhister	budhists,buddhists,
listor	lists,
personal	staff,
förödande	devastating,
amerikanen	american,
amerikaner	american,
irans	iran's,
förstnämnda	first-named,aforementioned,
aborter	abortions,
infektioner	infections,
aston	aston,
startat	started,
medlemmar	members,
downs	down,
stimulerar	stimulates,stimulating,
omgivning	surroundings,ambient,surrounding,
isen	the ice,
lärjungar	disciples,
huvudrollen	the main role,
inledde	launched,
tillvaron	existence,the subsistence,
sida	page,side,
överraskande	surprisingly,
bröllopet	the wedding,wedding,
side	side,
kammaren	chamber,the chamber,
centralt	centrally,
huvudstaden	capital,
liga	compatible,
päls	fur,
enorm	huge,
medier	medias,
milan	milan,
aids	aids,
håret	the hair,
kiev	kiev,
uppsala	uppsala,
hänvisa	reference,
talet	rate,
ihop	up,together,
talen	rate,
återfanns	was rediscovered,found,can be found,
venezuela	venezuela,
bestod	was,
normer	norms,standards,
stöds	supported,stood,
nomineringar	nominations,
folkvalda	elected,popularly elected,
faktum	fact,
iso	iso,
reinfeldt	reinfeldt,
representant	representative,
uppbyggt	structured,
starta	start,launch,
gå	go,
nätet	net,
jordanien	jordan,
arrangeras	(is) arranged,
skalvet	quake,
leddes	was led,
återkomst	return,
objektet	object,
föreslagit	suggested,
girls	girls,
vikingatiden	the viking age,
förbi	past the,
objekten	objects,the objects,
hollywood	hollywood,
någonstans	somewhere,nowhere,
åskådare	audience; viewer,
medeltiden	middle ages,
besegrades	defeated,
skaffade	aquired,
grönwall	grönwall,
symptom	symptom,
hundar	dogs,
formell	formal,
kontrast	contrast,
antarktis	antarctica,antarctic,
regissören	director,
härkomst	provenance,
parter	party,sides,
troligtvis	probably,
palace	palace,
stadsdelen	the district,district,
mina	my,
modern	modern,
självständiga	independent,sjalvstandiga,
brittiske	british,
självständigt	independently,independant,
triangel	triangle,
tecken	characters,signs,
lämnas	left,
lämnat	left,
skildringar	description,scenes,
tidiga	early,
monetära	monetary,
muskler	muscles,
förefaller	appear,
tidigt	early,at an early stage,
tål	is resistant to,stand,can take,
blue	blue,
bildas	formed,
tåg	rail,
bildat	formed,
mario	mario,
luthers	luthers,
marie	marie,
typ	type,
diskuterats	been discussed,
maria	maria,
don	don,
dom	judgement,conviction,
materiella	material,
talanger	talents,
spontant	spontaneously,
slipknot	slipknot,
vänta	(have to) wait; expect,wait,
följande	the following,
dos	dosage,
dop	baptismal,
kristen	christian,
långvariga	long,
koppla	coupling,
införde	enforced,introduced,
västeuropa	western europe,
kronprins	crown prince,
liza	liza,
droger	drugs,
nevada	nevada,
odling	cultivation,
krönika	chronicle,
förutsätter	assume,assumes,
folke	folke,
helhet	entirety,
monica	monica,
stycke	piece,piece; part; section,
kollapsade	collapsed,
stop	stop,
stol	seat,
strategiska	strategic,
mönster	marks,
earl	earl,
bar	bar,
bas	base,
existerar	exists,
skrivas	written,printed,
existerat	existed,
noga	carefully,
bad	bath,
fokus	focus,
liggande	placed,overhead,lie,
gärningar	yarn penetrations,deeds,
playstation	playstation,
zonen	zone,
zoner	zones,
gunnar	gunnar,
vända	turn,
dittills	thus far,so far,
vände	reversed,turned,
öppnade	opening,
inledningsvis	initially,in the beginning,by way of introduction,
naturligtvis	off course,naturally,
skrift	book,writing,
sorts	variety,
göta	göta,
omkringliggande	surrounding,neighbouring,
smguld	sm gold,
artikel	article,
armeniska	armenian,
nationalister	nationalists,
harvard	harvard,
kämpa	fight,
motto	motto,
regelbundet	regularly,
isotoper	isotopes,
regering	the government,
näringslivet	industrial life,
fördraget	the treaty,treaty,
fördragen	treaties,the compacts,
ernst	ernst,
upptäcker	discoveries,
kopplingen	the connection,
mellanrum	gap,
nationalförsamlingen	national assembly,
synsättet	view,
avsikt	intention,intends,
olsson	olsson,
varmt	hot,warm,
basis	basis,
sidan	page,
blodkroppar	blood cells,corpuscle,
cyrus	cyrus,
ting	things,
tina	defrost,
tillämpa	administer,implement,
idol	idol,
minoriteten	minority,
betydelsefull	significant,
igång	start,start up,
provinsen	province,
provinser	provinces,
sällskapshundar	pet dogs,
namnen	the names,
mindre	smaller,less,
etniskt	ethnic,
blåvitt	blåvitt,bluewhite,blue and white,
etniska	ethnic,
pornografi	pornography,
paradiset	the paradise,paradise,
förgäves	in vain,
albaner	albanians,
kvinnor	female,women,
ip	ip,
sushi	sushi,
it	it,
ii	(ii),
cant	cant,
dokument	files,document,documents,
il	il,
sommar	summer,
indonesiska	indonesian,
utgåva	edition,issue,
stoppa	stop,
konkurrensen	competitive,
vänstern	the left wing,left party,
make	husband,
producerats	produced,produced (by),
bella	bella,
kommunistpartiets	communist party,the communist party,
roland	roland,
därmed	consequently,therefore,
makt	power,
benämningar	names,
atmosfären	atmosphere,
försvarets	forsvarets,
skickades	sent,
nicklas	niclas,
akademiska	academical,academic,
protesterna	the protests,
nedan	below,hereinafter referred to as,
sydamerika	south america,
fuglesang	fuglesang,
glädje	joy,
dåvarande	then,
värmland	varmland,värmland,
roma	roma,
viktiga	important,
grannländer	neighbors,neighboring countries,neighboring lander,
just	currently,just,
diameter	diameter,
jämför	compare,
universitet	university,
psykos	psychosis,
bollen	ball,
västeuropeiska	western european,
viktigt	important,
human	human,
anders	anders,
beskriver	describes,
premiärminister	prime minister,
fysiker	physicist,
hävdar	states,maintain,
bokstäver	letters,
troligt	likely,
hävdat	claimed,
självstyrande	self-governing,
strax	soon,just,
royal	royal,
julen	julien,christmas,
memoarer	memoirs,
jules	jules,
friedrich	friedrich,
borgen	the castle,
komintern	comintern,
språkets	language,
arkitekturen	architecture,
behövde	did,needed,
rättegång	trial,
särdrag	feature,features,
följaktligen	consequently,
tittar	looking; viewing; viewer,viewing,
författningen	constitution,
gustaf	gustaf,
trafikeras	served,
trafikerar	traffic,
världsdel	continent,
sjöfarten	maritime transport,shipping,
medborgarskap	citizenship,
kommunerna	kommunera,
släkting	relative,
intensiv	intensity,
juryns	the jury's,jury,
syrien	syria,
kemiska	chemical,
vattnet	water,the water,
kontinent	continent,
dead	dead,
uppmärksammades	attention,
jupiter	jupiter,
befann	found,located,
kemiskt	chemically,
dominerade	dominated,
tappar	drop,lose,
statistik	statistics,
oralsex	oral sex,
hudfärg	color,skin color,
miljöproblem	environmental problem,
normal	normal,
arthur	arthur,
däggdjuren	the mammals,
säsongerna	seasons,sason organize,
filmatiserats	been filmed,screened,
benämns	designated,is mentioned,
mynt	coin,
angrepp	attack,
burj	burj,
versioner	versions,
bolt	bolt,
härstamma	originate,stem,
burr	burr,
förkortas	reduced,
super	super,
irländska	irish,
fördelen	advantage,
ljungström	ljungstrom,ljungström,
avgör	decides,avor,
därutöver	in addition,
maskiner	machines,
omröstning	vote,
tolkats	interpretation,
tillverkar	producing,
magazine	magazine,
ishockey	ice hockey,
grenen	branch,
förknippade	associated,
äktenskap	marriage,
psykisk	mental,
romantiska	romantic,
français	francais,public,
guide	guide,
jens	jens,
orsak	reason,
utbildning	eduction,
amsterdam	amsterdam,
havsnivån	sea level,
fastlandet	mainland,
estniska	estonian,
tennis	tennis,
bolivia	bolivia,
märke	badge,label,
hyllade	celebrated,acclaimed,
form	form,
norrlands	northern sweden's,norrland,
batman	batman,
ford	ford,
berg	mountain(-s),mountain,
japansk	japansk,japanese,
bero	due,
bättre	better,
byggde	built,
definierade	defined,
tempel	temple,
spelade	played,
positiv	positive,
flickvän	girlfriend,
åriga	year,
regeringen	government,
båten	vessel,boat,
skelett	skeleton,
beteckningen	the label,designation.........,designation,
frihetliga	libertarian,
försörjde	living,
handelspartner	trading partner,
tosh	tosh,
kanske	may,
mänsklighetens	humanity's,
tämligen	rather,tamil again,
vista	vista,
handen	hand,
handel	commercial,
kunnat	could have been,
betala	pay,
digital	digital,
betalt	charge,
marxism	marxism,
kungamakten	monarchy,
överenskommelse	deal,
frodo	frodo,
accepterade	accepted,
lokal	local,
engagemang	commitment,
riktad	directed,
ökande	increasing,rising,
ansökte	applied,
prov	test,
riktat	riktag,
riktas	target,
fattas	taken,
milt	mild,
armar	arms,
bomben	the bomb,
telefon	telephone,
tredje	third,
manager	manager,
bomber	bombs,
vikingarna	the vikings,
marissa	marissa,
dä	the elder,
då	when,
avbrott	breaks,
uppdelning	division,
petersburg	petersburg,
belgiens	belgium's,
din	yours,your,
fackföreningar	unions,
dig	up,
trenden	the trend,
afrikansk	african,
höjdes	increased,
dit	there,
spets	edge; top,tip,point,
bulgarien	bulgaria,
ville	wanted (to),wanted,
malmö	malmo,
diskografi	discography,
villa	house,
slagit	held,beaten,
reklamen	the commercial,commercial; ad; advertisment,advertising,
invandringen	immigration,
rymden	space,
hästen	the horse,
bakom	behind,
afghanistan	afghanistan,
viktig	important,
södra	southern,south,
föredrog	prefered,
bibliotek	library,
lönneberga	lönneberga,
somalia	somalia,
international	international,
madagaskar	madagascar,
avsluta	exit,
nationalismen	nationalism,
högkvarter	headquarters,head quarter,
avsaknad	absence,
kommun	local,
beskrivits	described,
boy	boy,
diagnoser	diagnoses,
bor	lives,
gyllene	golden,
partnern	partner,the partner,
mängder	amounts,amount,
extrem	extreme,
bob	bob,
diagnosen	diagnosis,
departement	departement,
sporter	sports,
enorma	enormous,
utövar	exercise,
utövas	exercised,
asiatiska	asian,
sporten	sport,port,
religionsfrihet	freedom of religion,
östasien	east asia,
platån	sycamore,
franco	franco,
hemmaarena	home ground,home field,
tennisspelare	tennis player,
socialister	socialists,
maya	maya,
peru	peru,
kristian	kristian,
förbjöds	banned,
detaljer	details,
avsattes	deposited,
ögon	eyes,
kemisk	chemical,
fartyget	ship; vessel,
fly	escape,
hända	may,provide,
hände	happened,
tokyo	tokyo,
mästarna	champions,
soul	soul,
träffades	met,was met,
vittnen	witnesses,
akademien	riksdagens,
präglade	characterized,
anslutna	affiliated,connected,
bristande	wanting,lack,
sökt	pending,searched,
hiroshima	hiroshima,
crazy	crazy,
kenneth	kenneth,
uruguay	uruguay,
winston	winston,
agent	agent,
skadades	was wounded,damaged,
council	council,
dennis	dennis,
kunglig	royal,
pink	piddle,
diskuterades	discussed,
oslo	oslo,
engelsmännen	the british,
varor	products,
ekonomiska	economic,
till	to,
gitarrist	guitarist,
nya	new,severe,
nye	new,
överensstämmer	agree,
fotboll	football,
läkare	doctor,
maj	may,
upphört	left the association,end,
man	is,
asien	asia,
johnson	johnson,
sådana	such,
eng	eng.,
q	q,
tala	speak,
basket	basketball,
romantiken	romance,romanticism,
nå	reach,
sådant	such,
lsd	lsd,
bussar	bus,
bevisa	prove,
alfabetet	alphabet,
städerna	city ​​limits,
sällsynta	rare,
protestantiska	protestant,protestantic,
lyrik	poetry,
motståndet	the resistence,
verksam	effective,
juryn	the selection panel,jury,
sekter	sects,
inkomster	revenue,
äkta	genuine,married,authentic,
nazisterna	nazis,
policy	policy,
main	main,
texas	texas,
lägst	lowest,lowermost,
steget	step,
kräver	requires,
janeiro	janeiro,
domstolar	courts,
mattis	mattis,
sibirien	siberia,
leds	passed,
färg	colors,colour,
leda	lead,
ledd	led,
föremål	object,subject,
tysklands	germanys,
guevara	guevara,
latin	latin,
tacitus	tacitus,
sökte	searched,
söner	sons,
vattendrag	watercourse,
avkomma	offspring,
girl	girl,
dianno	di'anno,
saudiarabien	saudi arabia,
enastående	outstanding,
håkansson	hakansson,
avrättningar	execution,executions,
områdena	the areas,areas,
tronföljare	heir,successor,
kattdjur	cat,
valdes	representatives',selected,chosen; elected,
ansiktet	face,
monster	monsters,
romani	romani,roma,
konstnär	artist,
chiles	chiles,
oro	anxiety,worry,
dubbla	double,
california	california,
miley	miley,
brooke	brooke,
befolkningens	population's,population,
ord	word,
tunnelbanan	subway; tube; underground,metro,
keith	keith,
verkade	were active, worked, was active,
gott	good,
upplevde	felt,
preventivmedel	contraceptives,preventivedel,
självmord	self-killing,
rankningar	ranking,
vision	vision,
stängdes	closed,
egentligen	actual,really,
föreställningen	the idea,the concept,show,
grupperna	groups,
intryck	appearance,
uttalanden	statements,
här	this; here,is,
rachel	rachel,
folklig	folk,
fast	solid,though; although; fixed; permanent,
grundämnet	the element,
missnöje	dissatisfaction,
visar	is,shows,
alfred	alfred,
grundämnen	elements,
individ	individual,
örebro	Örebro,
bobo	bobo,
anus	ass,
köpenhamns	copenhagen's,
fysiska	physical,
fysiskt	physically,physical,
löstes	solved,dissolved,
drevs	concentrated,was driven,
beslutet	the decision,
passade	suiting,suited,
fiender	enemies,
medlemmarna	members,the members,
lugn	calm,
jordytan	earth's surface,
fordon	vehicle/-s,vehicle,
inträde	entry,
marklund	marklund,
jämlikhet	equality,
stadsdelar	districts,city districts,neighborhoods,
större	greater,
formerna	forms,
tänder	teeth,
orsakerna	the causes,
kevin	kevin,
adeln	nobility,
nikola	nikola,
politiska	politic,political,
förälskad	in love,
menas	means,
skulptur	sculpture,
centralbanken	centralbank,central bank,
potential	potential,
performance	performance,
magnetiska	magnetic,
isolerad	isolation,isolated,
hertig	duke,
dagbladet	daily paper,dagbladet,
halvan	the half,
politisk	political,
teoretiskt	theoretic,theoretical,
mordet	the murder,murder,
beskrivit	described,
queens	queen,
över	over,
döden	death,
otaliga	countless,
lojalitet	loyalty,
drottning	queen,
grammatik	grammar,
österut	eastwards,
kontrolleras	controlled,
kontrollerar	controlling,
adolfs	adolf,
uranus	uranus,
regioner	regions,
generalsekreterare	the secretary-general,secretary general,
samlingsalbum	compilations,
helig	holy,
passande	suitable,
historien	history,
statsmakten	the government,
karolinska	caroline,
ges	given,be given,
ger	gives,
raser	races,
kulturellt	culturally,
konsolen	bracket,
motsvarande	corresponding to,
skådespelare	actor,
ramadan	ramadan,
personliga	personal,
katla	katla (fictive dragon in the classic "bröderna lejonhjärta"),
vintergatan	milky way,
firade	celebrated,
ledaren	leader,conductor,
rasen	breed,the race,
himmlers	himmlers,himmler,
försörjning	sustention,supply,
tillåta	allowing,
statistiska	statistical,
förenta	united,
spridda	spread,scattered,
världskrigen	the world wars,
europacupen	european cup,
london	london,
tolfte	twelth,twelfth,
relativt	relatively,
sämre	poor,samre,
sekulära	secular,
hittar	found,
fokuserar	focuses,
toppade	topped,
relativa	relative,
sean	sean,
slöt	joined (in peace),closed,
menat	meant,
menar	mean,
kandidater	candidates,
försvarsmakten	national defence,
visades	was,showed,
vanns	was won,
människan	the human,
söndagen	sunday,
personligt	private,
världskriget	world war,
gaga	gaga,
människas	human,
landets	its,
tsaren	the czar,czar,the tsar,
august	august,
 °c	celsius,
ju	the,
tur	tour,luck,
forskaren	researcher,
åker	treats,field; going,
timme	hour,
tum	inch,inches,
signaler	signals,
lexikon	lexicon,
ja	yes,
rugby	american fotboll,rugby,
ån	on,from,
utvalda	selected,selected; chosen,
tour	tour,
åt	to,for,
ås	ridge,
år	the year,
vätska	fluid,liquid,
naturresurser	natural resources,
jobb	job,
monarki	monarchy,
väst	west,the west,
cancer	cancer,
syntes	synthesis,
grundare	founder,
territorium	state,
mätningar	measurements,
ryggen	the back,
överföra	transmit,
bildats	had formed,created,
kirsten	kirsten,
industrin	industry,
västliga	western,
mars	march,
överförs	transfered,
plötsligt	sudden,
mary	mary,
flaggan	flag,
cobain	cobain,
avskaffa	abolish,
bmi	bmi,
klädsel	cover,
meningen	sense,
skriver	write,
sound	sound,
avsåg	mean,
dragit	dragged,preferred,
uppstod	was,
insåg	realized,
nionde	ninth,
sahara	sahara,
intressanta	interesting,
uppmanade	urged,encouraged,
liknande	similiar,similar,
uppfyller	fulfills,
hålls	is held,
par	pair,
upplagor	issues,
jesu	jesu,jesus,
edwin	edwin,
lava	lava,
hålla	hold,keep,
röka	smoking,
pan	pan,
samt	also,
hösten	fall,
running	running,
kuba	cubans,
teknisk	technical,
lösningar	solutions,
markus	marcus,
bang	bang,
wahlgren	wahlgren,
identifiera	identification,
gates	gates,
münchen	munchen,munich,
bebyggelse	habitation,
privatliv	private,
reaktionen	reaction,the reaction,
dinosaurierna	dinasaurs,
skapelse	creation,
vilja	will,like,
byggnad	building,
våld	violence,force,
jakten	the hunt,hunt,
ideologiskt	ideologically,ideological,
grannländerna	neighbors,
bowie	bowie,
avskaffandet	abolition,abolishment,
programledare	host,
bestämde	determined,chose,
motverka	prevent,counter,
trä	tra,
möter	meets,
schwarzenegger	schwarzenegger,
underarten	subspecies,sub species,
mor	mother,
haft	had,
prägel	character,mark,
mot	against,
temperatur	temperature,
mon	mon,
baltiska	baltic,
kollektiv	public,
mod	courage,mod,
christina	christina,
adams	adams,
födda	born,
började	began,
jordbävningar	earthquakes,
klubbarna	the clubs,
mänsklig	human,
sågs	seen,
göras	made,be made through,
grannar	neighbours,
kategorisveriges	category sweden,
joan	joan,
feodala	feudal,
konspirationsteorier	conspiracy theories,
förs	out,rapids,
jordbruket	the agriculture,
lotta	raffle,lotta,
fört	led,lead,
ställdes	prepared,
sudan	sudan,
föra	pre,
före	ahead (of), before,
ända	up,
demokratisk	democratic,
traditionell	conventional,
ände	of,end,
moderata	moderate,moderates,
vistas	live,present,
förlust	loss,
londons	london's,
inkomstkälla	source of income,was added to cold,
olof	olof,
tongivande	influential,
island	icelandic,
allians	alliance,
lands	on land,
lagarna	the laws,
retoriken	rhetoric,
auschwitz	auschwitz,
matematiska	mathematical,
arvid	arvid,
wilde	wilde,
einstein	einstein,
mark	ground, soil, territory,
jagar	hunts,hunting,
gravid	pregnant,
behandling	treatment,
varelse	creature,
emellanåt	once in a while,occasionally,
anfalla	attack,
fullständiga	full,
eget	own,
inletts	started,initiated,
utbredd	spread,
härifrån	here,
egen	own,
tävlingen	competition,contest,
exemplar	copies,
bibliografi	bibliography,
manuel	manuel,manual,
verkliga	fair,
kröntes	crowned,
humanismen	humanism,
håkan	håkan,
följde	followed,
manliga	male,
öns	island's,
prestigefyllda	prestigious,
skriven	written,
palats	palaces,palace,
sångerska	songstress,singer,
videon	the video,video,
film	film,
again	again,
genrer	genres,
effekt	effect,
istanbul	istanbul,
muren	wall,
produktiv	productive,
stannade	stayed,
spåret	groove,
genren	genre,
faktorer	factors,
däremot	however,
ordna	arranging,arrange,
profet	prophet,
ungarna	the young,
förändrade	altered,
rykten	rumors,
ledning	conduit,guidance,
henriks	henry,
kyros	cyrus,
chris	chris,
medicinska	medicinal,medical,
araberna	arabs,
palestinska	palestinian,
uppfostran	upbringing,
u	u,
medicinskt	medical,
kuwait	kuwait,
snabbaste	rapid,fastest,
begå	commit,
resolution	resolution,
åtskilda	separated,segregated,separate,
mellanöstern	middle,the middle east,
vila	rest,
socialismen	socialism,
inspirerat	inspired,
vill	to,
hindrar	stop; prevent,
ingripande	negative,intervention,
inspirerad	inspired,
levern	the liver,liver,
zink	zinc,
symbolen	the symbol,
symboler	symbols,
fortsatt	further,
seriens	series,
kasta	throw,
avhandling	thesis,
handlade	was (about); traded,was,
israeliska	israeli,isrealic,
fall	where,
ramen	frame,
stödja	support,
ramel	ramel,
kulminerade	culminated,
ansvarig	charge,
miljoner	one million,
båtar	boats,
bröderna	brothers,
suttit	been,sat,
ockuperades	occupied,
massor	(in) masses,tons,
växthuseffekten	the greenhouse effect,greenhouse effect,
intressant	interestingly,of interest,
material	material,materials,
abc	abc,
danmark	denmark,
abu	abu,
lärare	teacher,
långhårig	rough,long haired,long-haired,
närhet	close,proximity,
vald	elected,
jonas	jonas,
kandidat	candidate,
benen	legs,
valt	chosen,selected,
sångare	singer,
historiker	historians,
jackie	jackie,
tillkännagav	announced,
sjukhuset	hospital,
enat	united,
rösterna	votes,
författaren	the author,author,
hyllning	tribute; homage,
eye	eye,
medlem	member,
torrt	dry,
innebar	was; meant; entailed,
utmärkelser	awards,
torra	dry,
landet	the country,
människa	man,
leonard	leonard,
koma	coma,
brist	non,lack,
udda	odd,
berätta	tell,
vladimir	vladimir,
der	where,
des	des,
det	it,
roosevelt	roosevelt,
lindgren	lindgren,
den	it,
lagerlöf	lagerlöf,
befintliga	current,existing,
samtliga	all,
hastigt	fast,
latinets	the latin's,
sovjetunionens	soviet union,
betoning	stress,
samhälle	society,
medförde	brought,led,
sträng	string,strang,
robinson	robinson,
protein	protein,
makten	power,
hämta	retrieve,
stil	type,
psykotiska	psychotic,
georgien	georgia,
stig	stig,
verkligheten	real,reality,
rapport	report,
undervisningen	teaching,the education,
vikten	importance,weight,
makter	powers,
hoppade	jumped,
avtalet	agreement,
pettersson	pettersson,
laboratorium	laboratory,
ännu	yet,
ligger	lies,
vatten	water,
rastafarianer	the rastafarian,rastafarians,
rockgrupper	rock groups,rock group,
paz	paz,
konservatismen	conservatism,
civila	civil,
bernadotte	bernadotte,
uppgav	said,
officiella	official,
fältet	the field,field,
förmågan	the ability,
göra	do,do; doing,
mörkt	dark,
tvåa	second,
baltikum	the baltics,baltics,
mörka	dark,
görs	made,is made to,
officiellt	official,
människans	human,
längden	lenght,
diskussion	discussion,
wilhelm	wilhelm,
edmund	edmund,
inbördeskriget	civil war; civil war,
epok	epoch,
odlade	cultured,
saknades	missing,
trossamfund	religious community,faith community,
suverän	terrific,supreme,sovereign,
good	good,
träffar	meets,hits,
planerna	plans,
fängelse	prison,
sexuellt	sexual,
oxford	oxford,
skrifterna	scriptures,
association	association,
porto	postage,
robbie	bobbie,robbie,
kungarna	the kings,kings,
inleder	start,
haile	haile,
mental	mental,
house	house,
energy	energy,
hard	hard,
byggs	building,under construction,
förenade	united,
energi	energy,
sanningen	truth,the truth,
tomt	blank,
×	x,
infrastrukturen	infrastructure,the infrastructure,
ölet	the beer,
forskning	research,
perro	perro,
förföljelser	persecution,persecutions,
fullständig	complete,
konflikt	conflict,
bränslen	fuel,fuels,
lawrence	lawrence,
strömning	strom accession,flow,
eventuella	any,
blekinge	blekinge,
uralbergen	the ural mountains,
eventuellt	possibly,eventually,
viken	gulf,
helsingör	helsingor,elsinore,
inflationen	inflation,
legender	legends,
utöver	addition,
harris	harris,
styre	rule,
legenden	legend,
ensam	alone,
styra	controlling,
top	top,
sjunkande	decreasing,
säkerhetsråd	security council,
snarast	rather,
carter	carter,
lidande	sufferer,
kom	came,
kol	coal; charcoal,
lördagen	saturday,
observationer	observations,
förhindrar	prevents,
kategoriasiens	category of asia,
costa	costa,
kardinal	cardinal,
järnvägar	rail,railways,
triangeln	triangle,
part	party,
domstolen	court,
början	top,
matteusevangeliet	book of matthew,
följden	the cause,
fattiga	poor,
knapp	scarce,bare,
proteinerna	the proteins,
dogs	dogs,
personens	the persons,
århundraden	centuries,
hellström	hellström,hellstrom,
baháí	baha'i,
avtar	declines,decreases,
självständig	independant,
följder	impact,consequences,
lyssnar	listens,
lägret	the camp,
försökte	try,tried to,
bränsle	fuel,
gjord	made,
flertalet	majority; plurality,several,
gjort	created,
mountain	mountain,
hundratals	hundreds of,hundreds,
mussolini	mussolini,
infrastruktur	infrastructure,
caesar	caesar,
genast	at once,immediately,
inkomsterna	the incomes,revenue,
hölls	was,
lettland	latvia,
varifrån	from where; wherefrom,
patterson	patterson,
krafter	forces,
gillade	liked,approved; liked,
niclas	niclas,
kraften	power,
utbrott	outbreak,outbreaks,
samtidigt	while,simultaneous,
organiserade	organized,
högt	high,
km	km,kilometers,
kl	at,o'clock,
kr	kronas,
höga	high,
organisk	organic,
thomas	thomas,
kvalitet	quality,kvalilet,
bergman	bergman,
relation	ratio,relation,
utveckla	developing,
fina	beautiful,fine,
nämns	mentioned,
antagit	adopted,
konto	account,
undre	lower,
wallenberg	wallenberg,
medverka	take part,participate,
världens	the world's,the world,the worlds,
tionde	tenth,
förbudet	ban,
avseende	regard,for,
toronto	toronto,
nationalpark	national park,
notation	notation,
beslutar	decides,
vänskap	friendship,
express	express,
beslutat	resolved,
förklarat	explained,declare,
typiska	typical,
förklarar	explain,explains,
gamla	old,
husen	housing,
wallander	wallander,
gamle	old,
uttrycket	the expression,expression,
uttrycker	express,expressing,express (-es),
flykt	escape,
huset	the house,
somrar	summers,
§ 	s,
suveränitet	sovereignty,
rollfigur	character,
godkännas	be approved,approved,pass on,
höglandet	highlands,
rovdjur	predator,
fans	fans,
landsbygden	rural,
champagne	champagne,
romarriket	the roman empire,
professionella	professional,
framförs	is presented,
framfört	expressed,presented,
rörelserna	the movements,movement,
framföra	express,
skivorna	the records,plates,
marilyn	marilyn,
musklerna	muscles,
statligt	state,governmental,
vuxit	grown,
restaurang	restaurang,restaurant,
baltimore	baltimore,
globala	global,
kroatiens	croatia's,croatias,
förklaring	statement,
folkmord	genocide,
karaktären	character,
andas	breath,breathes,
karaktärer	characters,
således	hence,thus,
tennessee	tennessee,
immunförsvar	immune defense,
behöll	kept,retained,
försäljningen	gush sales,
lyfta	lift,
våningar	floors,storeys,
laos	laos,
fördrevs	ford described,
inför	before,
popularitet	popularity,
gav	gave,
effektiva	effective,
gas	gas,
vana	familiar,used,
kalmar	kalmar,
vann	won,
detsamma	the same,same,
bild	picture,image,
motorväg	freeway,highway,
åtalades	was prosecuted,
spridning	proliferation,
döptes	renamed,
portugal	portugal,
arenan	arena,
elektronik	electronics,
påbörjade	started,
monroe	monroe - it's a persons name,
rederiet	the shipping company,the company,shipping company,
dödat	killed,
granska	exam,
sjuk	ill,disease,
dödar	kill,kills,
tänkt	supposed; intended,intended,
administrationen	administration,
dödad	killed,
tyder	indicates,
sittande	fitting,
övertogs	were taken,
skotska	scottish,
syd	south,
konstnärliga	artistic,
syn	sight,view,
jerusalems	jerusalem's,
moment	step,
kallades	called,
kraftig	strong,
nämnde	mentioned,said,
nämnda	said,
kungariket	kingdom,
noll	zero,
kapitel	chapter,
albanien	albania,
jorderosion	earth erosion,soil erosion,
värme	heat,thermal,
skott	bulkheads,round,
albanska	albanian,
norrland	northern,
dikter	poems,
kommunister	communists,
juventus	juventus,
halvt	half,
ande	of,
verkställande	executive,
passerar	passes,
struktur	structure,
senaste	last,
alternativt	alternatively,
analytiska	analytical,
alternativa	alternative,
tropisk	tropical,
sektion	section,
kubas	cuba,cuba's,
monarkin	monarchy,the monarchy,
dömd	sentenced,
administrativa	administration,administrative,
dubbelt	double,
bil	car,
teknik	technique,technology,technic,
big	big,
kejsaren	the emperor,
avlidna	diseased,the perished,
möttes	met,
bit	piece,
planeterna	planets,the planet's,
rené	rené,
princip	principle,principal,
möjlig	possible,
stränga	severe,
tillstånd	condition,
figurerna	figures,characters,
google	google,
identisk	identical,
egyptiska	egyptian,
studerar	study,studies,
cocacola	coca-cola,
lars	lars,
västergötland	västergötland,
flygplatser	airports,air ports,
måste	have to,must,
per	per,
pratar	talks,talking,
diplomatiska	diplomatic,
energin	the energy,energy,
lösningen	solution,
nordamerika	north america,
resande	travelers,
vasaloppet	vasaloppet,
påven	the pope,pope,
ockuperade	occupied,
britannica	britannica,
drama	drama,
värmestrålningen	heat radiation,
uppfattningar	opinions,perceptions,
fallit	fallen,fall,
jimmy	jimmy,
grammy	grammy,
styrelse	government; direction,board,
barcelonas	barcelona's,barcelona,
steven	steven,
ordnar	fix,decorations,arrange,
paret	pair,the couple,parathyroid,
ökningen	increase,the increase,
dalar	valleys,
turkiska	turkish,
medvetande	consciousness,awareness,
jaga	course,chase,
serie	comic; row; succession; serial,series,
konsul	consulting,consul,
bostäder	housing,
torsten	torsten,
oktober	october,
skillnaden	the difference,
ledningen	the lead,conduit,
mångfald	variety,
smycken	jewlery,jewellery,
sultanen	sultan,
planer	plans,
amfetamin	amphetamine,
skillnader	differences,
reggaen	reggae,the reggae,
jordbävningen	earthquake,
reidar	reidar,
titel	title,
expedition	expidition,
förbjudna	forbidden,prohibited,
hjärnans	brain,
tropiskt	tropical,
materia	materia,
eller	or,
voltaire	voltaire,
familjer	families,
årstiderna	the seasons,arstiderna,
familjen	the family,
makedonien	macedonia,
anser	believes,view,
tvserie	tv serial,
maos	mao,
lena	lena,
länders	countries',countries,
samla	collecting,collect,
mutationer	mutations,
nådde	reached,
ritualer	rituals,
regionala	regional,
sambandet	relation,
dramatiker	dramatists,
judisk	jewish,
sorg	grief,sad,
regionalt	regional,regionally,
flod	basin,
uppgår	is,shall amount,
jason	jason,
stänga	off,
stred	fought,
frankrike	france,
sigmund	sigmund,
stängt	closed,
intensivt	intensive,
privat	private,
lilla	small,
tillämpningar	situations,implementations,
medlemskap	membership,
betrakta	view; regard,view,
sydafrikanska	african,
sahlin	sahlin,
konsten	art,the art,
intensiva	intensive,
kollaps	collapse,
atlas	atlas,
graven	grave,
luleå	luleå,
kampanjen	campaign,
plikt	duty,
släppte	released,
tjänade	earning,earned,
utgjordes	make up,comprised; consisted,
svts	svt,svts,
tävlingar	competitions,
exemplet	example,
joel	joel,
samman	together,
slutade	ending,
månens	the moon's,
warszawa	warsaw,
endast	only,
joey	joey,
tunnlar	tunnels,
störtades	overthrew,was overthrown,
överhöghet	suzeranity,
utbredda	spread,
vanligaste	frequent,
påsken	easter,
earth	earth,
carlo	carlo,
depression	depression,
edison	edison,
går	is,
chicago	chicago,
tillkomst	established,
placering	position,placement,
börje	börje,borje,
och	and,
kyrka	church,
öar	islets,islands,
extremt	extremely,extreme angular,extreme,
ordförande	chairman,
börja	start,
extrema	extreme,
isländska	icelandic,
populäraste	rated,
störning	noise,high accession,
honom	him,
svårigheter	difficulties,
medeltid	medieval,
alaska	alaska,
lagförslag	bill,
miljard	billion,
honor	female,
existens	existence,
protokoll	protocol,
uppnår	achieve,
talare	speakers,speaker,
privata	private,
hennes	her,
når	when,
nås	reached,is reached,
filippinerna	filipinos,the philippines,
betraktas	considered,
betraktar	regard,sees,
ovan	above,
lima	lima,
somrarna	summers,
kinesisk	chinese,
skotsk	scottish,
chi	chi,
gruppspelet	group stage,group play,
fånga	capture,capturing,
söder	south,
nytta	good,from,
geografisk	spatial,
titanics	titanic's,titanic,
prinsen	prince,
ledamöterna	the commissioners,commisioners,the members,
förstå	understand,first,
bakterier	bacteria,
avsikten	purpose,
engels	engels,
ansvaret	responsibility,the responsiblity,
britney	britney,
f	f,
tunnel	tunnel,
gabriel	gabriel,
påbörjas	starts,begin,
arton	eighteen,
baserad	based,
kedja	chain,
kategorisvenska	category: swedish,
baseras	based,based on,
baserar	base,
baserat	based,
kyrkan	the church,
vissa	some,
fotosyntesen	photosynthesis,
titlar	titles,
mozarts	mozart's,
cecilia	cecilia,
fett	fat,
internationellt	international,internationally,
lanserade	introduced,launched,
internationella	international,
tjänst	tjanst,
vilhelm	vilhelm,
revs	described,was demolished,
böckerna	books,
riktig	real,
frac	fraction,
malta	malta,
föddes	born,
herrlandskamper	men's international contest,men's international contests,
brändes	burned,burnt,
spannmål	grain,
förbundskapten	manager,
klan	clan,
gammal	old,
terrier	terriers,terrier,
siv	siv,
finländska	finish,finnish,
rådhus	townhouses,town hall,courthouse,
dryck	beverage,drinks,
förekommit	occured,
registrerade	data,
olyckan	incident,the accident,
alltjämt	remains,
bilbo	bilbo,
omslaget	cover,
dy	younger,
halvklotet	hemisphere,
strid	conflict,fight,
le	le,
variationer	variations,
berget	mount,
föreställer	pictures,depicts,
tillägg	addition,
weber	weber,
dag	dag,day,
referenser	references,
spela	play,
dam	lady,
dan	dan,
avslöjar	reveals,
tillkommit	been,accured,
periodiska	periodic,
sammanhanget	connection,
installera	installing,
day	day,
kontinuerligt	continuous,
beslut	decision,
morris	morris,
newtons	newton,
spridningen	the spread,
warner	warner,
engelskspråkiga	english-speaking,
juridisk	legal,
krita	chalk,
humanism	humanism,
pitts	pitts,
kristiansson	kristiansen,
dokumentär	documentary,
inspirerade	inspired,
segern	the victory,victory,
programmet	program,the application,the program,
arbetskraft	labor,
fattigdomen	poverty,
nödvändiga	necessary,essential,
matt	matt,dull,
jerusalem	jerusalem,
mats	attention,
kärnan	core,
ren	deer,clean,
deras	their,
red	eds,
återta	retake,regain,
roterande	rotating,
webbplats	site,
franz	franz,
odlas	cultured,
arbetare	workers,
ronald	ronald,
längre	longer,
josé	jose,
efterträddes	succeeded,
medelhavsområdet	mediterranean,
farbror	uncle,
fotografier	photographs,
south	south,
liberaler	liberals,
stämmer	(if it's) true,is true,
pga	because of (short of "på grund av"),
uppger	states,state,
innehålla	contain,
levnadsstandarden	living standard,
omständigheter	circumstances,
leder	leads,leading (to),lead,
utlopp	outlet,
energikällor	energy resources,
drabbade	affected,
förklara	declaring,explain,
maidens	maidens,
leden	lines,the route,
palestina	palestine,
demonstrationer	demonstrations,
bundna	tied,bonded,
släktet	the genus,
stället	instead,
ställer	run (in election),
innehade	held,possessed,
firades	celebrated,was,
treenigheten	tinity,the trinity,trinity,
tätorter	cities,
sjögren	sjögren,
ledamöter	commissioners,
släkten	genera,
ambassad	embassy,
domaren	the judge,
matematisk	mathematical,
uteslutande	only,exclusively,
kvalificerade	qualifying,
mälaren	mälaren,
premiär	prime,premiere,
havs	at sea,
aristoteles	aristotle,
biologiska	biological,
operativsystem	operative systems,os,operating system,
följd	consequence,effect,
älgar	moose,
följa	following,follow,
basist	bassist,
uganda	uganda,
rådande	current,
följt	followed,
följs	followed,
låt	let,
mil	mil,
min	my,
fötter	feet,
tidningar	press,magazines,
mig	me,
mix	mix,
låg	low,
experter	experts,
besättningen	crew,
lån	loan,
konstverk	artwork,
kommunikationer	communications,
resurser	resources,
dinosaurier	dinosaurs,
varandras	each others,each other,
missionärer	missioners,missioner,missionaries,
resultaten	the results,
sedan	then,
sist	finally,
herman	herman,
liknade	looked like,similar,
stranden	shore,the beach,
upprustning	renovation,
irakkriget	iraq war,
republikanska	republican,
rörelsens	movement,
milano	milano,
deuterium	deuterium,
tidskrift	magazine,
capita	capita,
styrke	strength,
definiera	defining,
viktigaste	most important,
styrka	strength,
utgångspunkt	starting point,point of departure,
obelix	obelix,
text	text,
komplicerad	complicated,
existerande	current,
inhemsk	native,
ugglas	ugglas,
timmar	hours,
kurfursten	elector,
rumänska	romanian,
järnvägen	rail,
euroområdet	euro area,
satan	satan,
shahen	the shah,shah,
säker	items,
bryssel	brussels,
organiska	organic,
djurgården	djurgården,zoo,
influensavirus	flu virus,flue virus,
förändrades	changed,
buddhismen	buddhism,buddism,
överlägset	far,
förstår	understand,forstar,
regimen	regime,
studenterna	the students,
uppehåll	residence,pause,
richards	richards,
från	from,
vinsten	gain,
organ	agency,organ,
majoriteten	the majority,
lyckade	successful,
byggdes	was built,
ronaldo	ronaldo,
militärer	military,
krävdes	were required,
national	national,
svenska	swedish,
eleonora	eleonora,
kapitalet	the capital,capital,
svenskt	swedish,
först	first,
bön	nests,prayer,
debutalbumet	debut album,
reform	reform,
redan	has already,
konverterade	converted,
raúl	raul,
bruno	bruno,
carlsson	carlsson,
avslutades	closed,ended; concluded,
bör	live,should,
terräng	off,
ordentligt	proper,properly,
översikt	overview,
koncept	concept,
industrialisering	industrialization,
uppskattade	estimated,appreciated,
hårdare	more severely,tougher,
säkerheten	the security,safety,
översättas	translated,translated (to),
viktigare	more important,
läsning	reading,
hämtade	taken,
buddhas	buddha's,buddhas,
empathy	empathy,
återförening	reunion,
litteratur	literature,litterature,
aktuellt	relevant,
kommunicerar	communicates,
aktuella	current,
kommendör	commandor,commander,
förekomst	presence,
sachsen	saxony,
dödsorsaken	cause of death,
befogenhet	authority,
utsågs	was,appointed,was appointed,
medicinsk	medical,
elektroner	electron,electrons,
västmakterna	western powers,
af	of,of (old swedish),
grupperingar	groupings,
slippa	avoid,
gaza	gaza,
igen	again,recognize,
define	define,
asteroider	asteroids,
genomsnittlig	average,
stationen	station,
stationer	stations,
orange	orange,
deep	deep,
an	an,
napoleon	napoleon,
augusti	august,
bruket	use,the use,
kraftiga	powerful,
stalin	stalin,
ar	is,
klassificera	classifying,classify,
betraktade	considered,watched,
externa	external,
kväve	nitrogen,
tagits	taken,
flyktingar	refugees,
verkligen	real,the reality,
fördrag	agreement,treaty,
partner	partner,
prosa	prose,
utom	out,
händelserna	the events,events,
administration	administration,
lämnade	did,left,
wolfgang	wolfgang,
blodtrycket	the blood pressure,blood pressure,
sångerna	song are,the songs,
fler	more,
hinduismen	hinduism,
kallad	called,
kontrollera	control,
framförallt	above all,in particular; above all,
helsingborgs	helsing borg,helsingborg's,
kallas	called,
kallar	calls,
center	center,
öde	fate,
seth	seth,
antonio	antonio,
sett	seen,
hoppas	hope,
omgångar	in turns; periods; mandates,cycles,
svensk	swedish,
undvika	avoid,
position	position,
deltar	participates,
innehåll	content,contents,
kontaktade	contacted,
folkrepubliken	people"s republic,
mystiska	mysiska,
wagner	wagner,
misshandel	assault,abuse,
grekiskans	greek,
flertal	several,majority group,
vanligt	normal,
kampf	kampf,
liverpools	liverpools,
reformer	reformers,
anhöriga	relatives,kin,
landområden	land,
streck	bar,
match	game,match,
förnuft	common sense,
uppträder	occur,performs,
dubai	dubai,
demens	dementia,
innehöll	contained a ban on,include,containing,
chrusjtjov	khrushchev,chrusjtjov,
likt	like,
journalist	journalist,
works	works,
uppträda	appear,
albumets	album,
starkaste	strongest,the strongest,
värt	worth,
etablerades	was established,
minsta	minimum,
est	est,
joachim	joachim,
löser	solves,
skildrar	depicts,describes,portrays,
gisslan	hostages,
internationalen	international,
definitionen	the definition,
nattetid	overnight,
definitioner	definitions,
starkare	strong,stronger,
leopold	leopold,
nordkorea	north korea,north koreans,
socker	sugar,
ärkebiskopen	archbishop,
glada	happy,
mäktigaste	powerful,
slutgiltiga	final,
andel	share,
anden	the holy spirit,spirit,
folkräkningen	census,the census,
medverkar	contributes,contribute,
alexanders	alexanders,alexander's,
förstärka	enhance,
socken	parish,
omgiven	surrounded,
tränger	forces forward,
världsliga	worldly,
ljusare	brighter,
föredrar	preferred,
vimmerby	vimmerby,
hatar	hate,
ridge	ridge,
densamma	same,
illuminati	illuminati,
kuben	the cube,
möjliggjorde	enabled,
flyg	airforce,
kärnor	cores,
klockan	clock,
brand	fire,
bröder	brothers,
ersättning	pay,replacement,remuneration,
flygvapnet	air force,the airforce,
kraft	force,power,
hinner	have time to,
nöjd	content,
vetenskap	science,
utrymme	space,
arbetsgivaren	employer,
individens	the individual's,
australiens	australia,australia's,
omfatta	cover,
kaffe	coffee,
minuter	minutes,
vänstra	left-hand,left,
hästens	horse's,
paraguay	paraguay,
tolkningen	interpretetation,interpretation,
omloppsbanor	orbits,orbit,
autism	autism,
vinner	wins,
manlig	male,
identitet	identity,
särskilda	specific,special,
proteinet	protein,the protein,
betonade	emphasized,
uppfattas	be perceived,are regarded,
försämrades	worsened,decreased,
uppfatta	apprehend,perceived,perceive,
sjön	sjon,lake,
astronomi	astronomy,
variation	diversity,variety,
koncentrationsläger	concentration,
akademisk	academic,
cirkel	circular,
särskilt	especially,
philips	philips,
fakta	facts,fact,
winnerbäck	winnerbäck,
svag	weak,
uppfattningen	comprehension,
framför	in front of,above,
förbundet	the union,association,
okänd	unknown,
brottslingar	criminals,
nederländerna	the netherlands,
båt	boat,
resor	travels,
påsk	easter,
arkitekt	architect,
antisemitiska	antisemetic,anti-semitic,antisemitic,
ozzy	ozzy,
anfallet	attack,
huvudstad	capital city,capital,
paris	paris,
tillväxten	growth,
under	under,
läge	mode,
svårare	answering machine,
pommern	pommern,pomerania,
ägande	ownership,
halsen	throat,
jack	jack,
invånare	inhabitants,
evert	everted,evert,
ovanstående	above,
tagit	taken,received,
school	school,
utmärks	are characterized,characterized,
utmärkt	excellently,
öppna	open,
plural	plural,
matematik	mathematic,mathematics,
verklig	real,
reklam	advertising,
parten	party,
markerar	selects,marks,
uppdelningen	partitioning; sectionalization; division; split (-ting),splitting,division,
bönderna	farmers,
manus	script,
läget	location,
indierna	indians,
läger	camp,
stridigheter	oppositions,strife,
aktivt	active,actively,
drivande	drive,
notera	note,
liberty	liberty,
aktiva	active,
sund	healthy,narrow,
kub	cube,
egyptens	egypts,
språken	languages,
zach	zach,
prata	talk,
flera	many,multiple,
medelhavsklimat	mediterranean climate,
utredning	study,investigation,
beck	beck,pitch,
parlamentariska	parliamentary,the parliamentary,
preparat	preparations,
studio	studio,
atombomberna	atomic bomb,
komplex	complex,komplex,
språket	language,
lagras	stored,
precis	just,
gällande	current,
upptäckter	discovery,
upptäcktes	discovered,(was) discovered,
julie	julie,
erektion	erection,
julia	julia,
övers	transl,translation,
nazistiska	nazi,
misslyckats	failed,
upptäckten	the discovery,
försvarsmakt	armed forces,
eftervärlden	posterity,
volym	volume,
klassas	classified,
vinst	win,
miniatyr|px|en	miniature,
konserterna	concerts,
västtyskland	västttyskland,west germany,
skicka	send,
behandlingar	treatments,
belägg	evidence,
övertala	persuade,
ludvig	louis,ludvig,
vagnar	carts,wagons,carriges,
världsarv	world heritage,
waterloo	waterloo,
igelkottens	hedgehog,
henri	henri,
mm	etc.,
arméns	the army's,
lukas	lukas,
antiken	the ancient world,antiquity,
ms	motor ship,
mr	herr,mr,
johanssons	johanssons,johansson,
avstå	non,refrain,
utgick	was deleted,
partiets	the party's,parties,
sträckan	distance,the distance,
utlöste	triggered,
persien	persia,
trädgård	garden,
florida	florida,
genomfördes	completed,was,
fröken	miss,
ena	one,
end	end,
smält	melted,
iiis	iii's,3's,
väpnade	armed,
ens	even,
gata	street,
elektriskt	electric,
elizabeth	elizabeth,
beskrev	depicted,described,
mest	most,
västvärlden	west,western world,
målet	target,
frågade	inquired,
 cm	centimeters,
kategorier	categories,
kubanska	cuban,
existera	exist,
arbetat	worked,
praxis	practice,
arbetar	works,
kejsare	emperor,
kampen	the struggle,the fight,fight,
arresterades	was arrested,
besittningar	holdings,possessions,
synonymt	synonymously,
frivillig	optional,
bär	berries,
brinner	on fire,
ursprungsbefolkningen	indigenous people,
imf	imf,
edith	edith,
nytt	new,
dött	died,
dem	those,
produktion	production,
upptagen	included,
livstid	life span,
ansvarar	charge,responsible,
alex	alex,
jämförelser	comparison,
detroit	detroit,
borrelia	borrelia,borreliosis,
storlek	size,
stadigt	steadily,stable,
gymnasium	high school,
dessförinnan	before,
träffade	met,
innehållande	containing,
raid	raid,
näst	second (to),
nio	nine,
medelålder	middle age,
god	good,
receptorer	receptors,
ammoniak	ammonia,
hemland	homeland,
riktning	direction,
danmarks	denmark's,
paulus	paulus,paul,
got	got,
behöva	need,
independence	independence,
snuset	snuff,the snuff,
icke	non,none,
värnplikt	military service,
free	free,
fred	peace,
statsöverhuvud	head of state,
undervisade	taught,
hört	heard,
inom	in,
drygt	good,
statsministern	prime minister,
studera	study,
tolerans	tolerance,
bredvid	beside,
vetenskapliga	scientific,
hjälpte	helped,
befolkade	inhabitated,populated,
vetenskapligt	scientific,
transporterar	carrying,
transporteras	transported,
säsong	season,
museet	the museum,museum,
museer	museums,musser,
nhl	nhl,
rikaste	the richest,
tillåts	allowed,
yngsta	youngest,
sexuella	sexual,
nyheten	news,
mercury	mercury,
toy	toy,
yngste	youngest,
punkten	the point,point,
konventionen	the convention,convention,
merkurius	mercury,
å	of the,
konventioner	conventions,
ton	tonne,
tom	tom,
uppkommit	generated,
tog	was,
fördes	sea were entered,
adjektiv	adjective,adjectives,
ifrågasatts	is questioned,
livealbum	live album,
skildes	was seperated,
rädsla	fear,
fördel	advantageously,
kulturarv	cultureheritage,
territoriella	territorial,
dramer	dramas,
slutsats	conclusion,
mjölk	milk,
uppmuntrade	encouragement,encouraged,
rad	line,range,
flyttades	moved,
tänka	thinking,
rak	linear,
somliga	some people,some,
störningar	disorders,
växer	growing,grows,
ras	race,ras,
övervikt	obesity,overweight,
motståndaren	adversary,
industriellt	industrial,
hittats	found,
kvällen	the evening,evening,
lanseringen	the release,launch,
användning	use,use; usage,
fartyg	vessel,ship,
industriella	industrial,
situationen	situation,the situation,
mekaniska	mechanical,
grundskolan	elementary school,
skepp	ship,
elektricitet	electricity,
fralagen	the fra law,
motsatt	opposite,
framgångsrik	successful,
motsats	contrary,
tanzania	tanzania,
metal	metal,
sjöar	lakes,parks,
inflytande	influence,power,
rikskansler	chancellor,
agnes	agnes,
utkanten	outskirts,
dyrare	expensive,
saga	story,
järnvägarna	the railways,railways,
queen	drottning,
gränserna	borders,the borders,
höjdpunkt	highlight,climax,high point,
sagt	said,
radie	radius,
erkänner	recognize,
claude	claude,
florens	florence,florens,
vinna	win,
resterande	remainder,
gods	goods,
holländska	dutch,
återstår	remains,
andras	others,
representerade	represented,represent,
kommunisterna	communists,
guatemala	guatemala,
gogh	gogh,
slags	kind,
ålder	age,alder,
stadskärnan	town/city,center,
ändras	be changed,
ändrar	changes,
ursäkt	excuse,apology,
ändrat	changed,modified,
lovat	promised,
utvisning	penalty,
kroppen	the body,
sakta	slowly,
ockuperat	occupied,
fördomar	prejudices,
utformade	formed,designed,
behålla	container,
mur	wall,
brinnande	burning,
antikens	the ancient's,ancient,
populär	popular,
slottet	castle,the castle,
finger	finger,finder,
förstås	course,
allra	very,
mun	mouth,
förhållande	ratio,(in) comparison (to),
ordnade	arranged,
betonar	stress,emphasize,
maniska	manic,
seden	the seed,custom,
inneburit	meant,resulted,
bildriksdagsval	image election,
kreativitet	creativity,
autonomi	autonomy,
anfall	attack,
verka	seem,appear,
lösningsmedel	solvent,
läggs	put before; submitted; put,lay,
allierades	allied's,allied,
begränsade	restricted,limiting,
förbränning	combustion,
viruset	virus,
lägga	put,lay,
katarina	katarina,
hitler	hitler,
solljus	sun light,sunlight,
skapades	generated,
rumänien	romania,
grundaren	the founder,founder,
strävhårig	hispid,wirehaired,
därefter	thereafter,
hastighet	speed,
diktatorn	the dictator,
homosexuell	homosexual,
skalan	scale,
öster	east,
modernare	mor modern,more modern,
anspråk	claims,
spritt	spread,
drömmar	dreams,
invasionen	invasion,the invasion,
älgen	moose,
petrus	petrus,
schizofreni	schizophrenia,
depp	depp,
claes	claes,
della	della,
nationer	nations,
viking	viking,
darwins	darwin,darwins,
därigenom	thereby,
vojvodskap	voivodships,
brott	breach,crime,
anlände	arrived,
nationen	the nation,
kartan	the map,
vanföreställningar	delusions,
varefter	whereafter,
ekonomin	economy,
väljs	selected,elect,
ernman	ernman,
återgick	returning,
pekar	points,pointer,pointing,
erhållit	acquired,received,
ökade	increased,
ersatte	substituting,replaced,
pekat	pointed,identified,
negativ	negative,
welsh	welsh,
hundra	hundred,
formatet	the format,
ersatts	replaced,(has been) replaced,
återvände	returning,
återvända	return,
uppsving	boost,
gudom	deity,
dylan	dylan,
charlie	charlie,
spelad	played,
svavel	sulfur,sulphur,
kemikalier	chemicals,
fattigare	poorer,
louisiana	louisiana,
jean	jean,
spelat	played,
spelas	played,
spelar	column,
mytologin	mythology,
kraftigt	heavily,
järn	iron,
torah	torah,
graden	rate,the degree,
europaparlamentet	european-parliament,the european parliament,european parliament,
grader	degrees,
engelskans	english,
utföras	performed,
kolväten	hydrocarbons,
kalifornien	california,
använt	used,
värnpliktiga	conscripted,inductees,
gavs	was,
eld	fire,
reglera	expell,controlling,
aktiv	active,
rätta	correct,come to grips; court; correct,
regionerna	regions,
enlighet	union,according,
 au	au,
tredjedelar	thirds,
donau	the danube,
ämnet	subject,
tillgänglig	provided,
protesterade	protested,
ämnen	agents,substances,
gift	married,
såväl	both,as well as,
ladda	load,
modersmål	native language,mother tongue,
bosnienhercegovina	bosnia-hercegovina,
specifik	specific,
tillåtna	allowed,
fotbollen	soccer,
gifter	marries,toxins,
lagstiftningen	law-making,
varianterna	variants,the diversities,
hanhon	he/she,male-female,
direkta	direct,
besöka	visit,
jennifer	jennifer,
malaysia	malaysia,
donald	donald,
besökt	visited,
saturnus	saturn,saturnus,
motsatsen	the opposite,
estetik	stetik,esthetics,
ultraviolett	ultraviolet,
totalt	complete,wholly,
användare	users,
icd	icd,
totala	total,
karaktäriseras	is charactarized,
elitserien	elite series,elitserien,
monoteism	monotheism,
ishockeyspelare	ice hockey player,hockey players,
tillbringar	spend,
män	males,men,
spelare	player,
hotellet	hotel,
titeln	the title,
tvingades	had,
systrar	sisters,
omgången	round,
plus	plus,
analytisk	analytical,
internationell	international,
tydliga	obvious,
genomslag	breakthrough,impact,
primitiva	primitive,
civil	civil,civilian,
menade	meant,
tydligt	obvious,
isberg	ice berg,iceberg,
sinne	mind,
oförmåga	failure,incapacity,
omger	surrounding,
lagt	added,
kjell	kjell,
sicilien	sicily,
anderson	anderson,
kronprinsessan	crown princess,
metabolism	metabolism,
wittenberg	wittenberg,
fadern	the father,
barrett	barett,barrett,
fängelsestraff	prison,
skulder	liabilities,debt,
finns	is,exist,there is,
eventuell	any,
fusionen	merger,the fusion,
säkerhet	safety; security,security,
amerikanerna	americans,
värvade	recruited,
araber	arabs,
behandla	treatment,
trio	trio,
bildt	bildt,
everest	everest,
bilda	form,
hamn	harbor,harbour,
kambodja	cambodians,
förbud	prohibiting,prohibition,
liberalism	liberalism,
tätorten	conurbation,
ni	you,
when	when,
nf	nf,
finna	found,
ny	new,
tio	ten,
tid	time,
nr	no,
höjer	rises,raise,raising,
nu	now,
picture	picture,
phoenix	phoenix,
sätts	is,turned (on),
miscellaneous	miscellaneous,
gäster	guests,
tunna	thin,
massakern	massacre,
sätta	insert,
väckte	aroused,
vietnam	vietnam,
cellens	the cell's,cell's,the cells,
rom	rom,
funktionerna	functions,the functions,
rob	rob,
dvärg	dwarf,
koreanska	korean,
tillkommer	will be,will be added,
fiktiv	fictitious,fictive,
mottagarens	the reciever,the receivers,
konstitutionell	constitutional,
tanke	in light of,
även	also,
underhållning	entertainment,
flytt	escaped,
krossa	crush,crushing,
metod	method,
inlärning	learning,
brother	brother,
christmas	christmas,
olyckor	accidents,
lever	liver,
länkar	links,
församling	congregation,
införandet	introduction,the introduction,
kategorirock	category rock,
colin	colin,
svartån	svartån (black stream),svartån,
uppgifterna	data,
ifråga	with regards to,
poesi	poetry,
agnosticism	agnosticism,
miniatyr	miniature,
ögat	eye,
cykel	bicycle,
månaderna	months,
angelina	angelina,
gräs	grass,
gravitation	gravitation,gravity,
kamp	struggle,fight,
vindkraftverk	wind power station,
enkla	simple,single,
metaller	metals,
eiffeltornet	the eiffel tower,
jord	earth,
dublin	dublin,
sina	their,
införts	introduced,
vägg	wall,
ankomst	arrival,
asterix	asterix,
tilltagande	increasing,
rafael	rafael,rafel,
luften	air,
etablera	erablera,establish,
trummor	drums,
bolaget	the company,
ungerska	hungarian,
russell	rusell,russell,
undan	away (from),escape,
utropades	was proclaimed,
samfundet	the communion,
abbas	abbas,
andy	andy,
kurder	kurds,
australian	australian,
turné	tour,
uppskattningar	estimates,
typerna	the types,types,
kär	in love,
övergå	transition,
palestinsk	palestinian,
årets	year,
efterhand	post,hindsight,
beroende	dependent on,depending,
styras	controlled,steered,
läkemedel	drugs,medicine,
musikaliska	musical,
rådgivare	advisor,
valla	wax,herd,
jude	dude,
allvarlig	serious,
domkyrka	cathedral,
humle	hop,
generell	general,
karibiska	caribbean,
anpassat	adapted,
uppväxt	growing up,
bönorna	bean,beans,
bära	carry,
dokumenterade	documented,
utdelades	awarded,
hemligt	secret,
annorlunda	different,otherwise,
hemliga	secret,
främja	promote,promoting,
swedish	swedish,
frivilligt	voluntary,
speglar	mirror,mirrors,
avrättning	execution,
frivilliga	volunteers,
andlig	spiritual,
stöter	run,
simning	swimming,
regeln	rule,
muslimerna	muslims,
inriktad	focused on,
tvserien	tv series,television program,
fascism	fascism,
sydliga	southern,
tvserier	tv-series,
flög	fly,
fenomen	phenomena,
leva	live,
utrikespolitiska	foreign policy,foreign political,
marknad	market,
riktar	target,
kroniska	chronic,
beror	is,
stridande	conflict,warring,
japanska	japanese,
representation	representation,
väntas	is expected,
väntar	waiting,expect,
faser	phases,
orter	varieties,locations,
kartor	maps,
bushs	bush's,bush,
orten	resort,the suburb,
födelse	date,
komplicerat	complex,complicated,
iberiska	iberian,
fasen	phase,
wallace	wallace,
försvinner	disappear,
klasser	classes,
spelarna	players,
försvaret	repository,the defense,
tjänstemän	officals,officials,
marleys	marley's,marley,
passar	suitable,suits,
hergé	herge,
femte	fifth,
hamilton	hamilton,
färgen	the color,
hotar	threatens,
opera	opera,operator,
snabb	instant,
futharkens	futhark,the futhark's,
viggo	viggo,
alternativ	alternative,
hotad	threatened,
färger	color,colors,
bildning	learning,form,
semifinal	semifinals,
förhandlingarna	negotiations,
stående	standing,
valuta	exchange,
rastafari	rastafarian,
amerikansk	u.s.,
åsikt	opinion,
tillhörighet	belonging,
behandlas	treated,
upprepade	repeated,
accepterad	acceptable,
stortorget	stortorget,
årliga	annual,
accepterar	accept,
accepterat	accepted,
kent	kent,
fortsättning	continuation,further accession,continued,
juldagen	christmas day,
etanol	ethanol,
nått	reached,
hjalmar	hjalmar,
gallien	gaul,
soundtrack	soundtrack,
arbetet	work,
händelse	event,
traditionen	the tradition,tradition,
motion	motion,exercise,
traditioner	traditions,the traditions,
place	place,
någonsin	ever,
politiken	policy,the politics,
arbeten	works,
blood	blood,
såldes	sold,
självbiografi	autobiography,
kontrollerade	controlled,
respekt	respect,
given	given,
ian	ian,
vågor	waves,
skjuten	shot,
sydafrika	south africa,
cullen	cullen,
bahamas	bahamas,
skjuter	shoots,
givet	granted,
folkmängden	population,
personlighetsstörningar	personality disorders,
webbplatser	webbsites,websites,
användandet	usage,use,
grund	in the context: "på grund" = because of,
montenegro	montenergo,montenegro,
alan	alan,
kallade	called,
hur	the,cage,
hus	house,a house,
webbplatsen	the website,site,
modellen	model,the model,
begravning	funeral,
marinen	navy,marines,
löfte	promise,
kontroll	control,
framställning	production,
landsting	county,county council,
bildades	founded,
hjärtat	heart,
rena	pure,
mottagare	recipient,
afrikanska	afrikanska,african,
tiotusentals	tens of thousands,
kromosomerna	the chromosomes,
kometer	comets,
rent	true,clean,
jordskorpan	the earth's crust,
världen	world,the world,
avstånd	distance,
förste	chief,
studion	the studio,
första	first,
fysikaliska	physical,
förhållandena	conditions,
gustavs	gustav,
kust	coastal,
periodvis	periodically,
stjärnornas	stellar,
knutna	tied,
fci	fci,
falla	fall,
fria	free,
staterna	usa,
täckt	covered,coated,
lisbet	lisbet,
elektromagnetisk	electromagnetic,
betydande	important,
stövare	beagle,hound,
täcka	cover,thank,
tron	faith,
ronaldinho	ronaldinho,
mänskligheten	humanity,manskligheten,
inåt	inwardly,
isolering	isolation,
tros	believed,
tror	think,
bandets	the bands,band,
gula	yellow,
guld	gold,
flydde	fled,
motivet	subject,
ovanligt	unusual,
gult	yellow,
iväg	away,off,
ovanliga	rare,
analys	analysis,
berättelser	tales,stories,
aktiviteten	the level of activity,activity,
grundandet	founding (of),founding,
tränaren	coach,the coach,trans breaker,
jazz	jazz,
administrativ	administrative,administration,
nedåt	down,downward,
väder	weather,
ansågs	was,
forsberg	forsberg,
beredd	prepared,
skivkontrakt	record deal,
dramat	drama,the drama,
joker	joker,
republika	republic,
osäkert	insecure,
satte	put together,
minnen	memories,
underlätta	ease,
tekniska	technical,
inspelningen	recording,
uppdraget	task; assignment,
stanley	stanley,
minnet	memory,
älg	moose,
freden	the peace,peace,
federal	federal,
utbud	range,
skett	happened,
hämtar	download,is,
återigen	yet again,aterigen,
intresserad	interested,
hämtat	collected,downloaded,
konstnären	artist,
antagligen	ligands presumably,probably,presumably,
konstnärer	artists,
bekämpa	prevent,fight,
ruiner	ruins,
dödade	killed,
myter	myths,
högre	higher,
summa	sum,total,
sydeuropa	southern europe,
region	region,
ordagrant	literal,
spindlar	spiders,
diskriminering	discrimination,
lenins	lenin,lenin's,
introducerades	introduced,
gjorde	did,
gjorda	done,
pakistan	pakistan,
utgåvor	editions,
regler	rules,
period	period,
pop	pop,
fransk	french,
werner	werner,
statens	state,
hävda	asserting,
poe	poe,
skånska	scanian dialect,scanian,skånska,
howard	howard,
förekomsten	presence,
dagarna	the days,day,
musikstil	music,
folket	the people,
invaderade	invaded,
andres	andres,other's,
hits	hits,
kapitulation	surrender,
tiger	tiger,silent,
övrig	other,
minister	minister,
kaos	chaos,
champions	campion,champions,
använder	using,
användes	was used,
riktade	targeted,
influenser	influence,influences,
cash	cash,
spreds	spread,disseminated,
fiende	enemy,
grundlagen	constitution,
odens	oden's,
universums	the universe's,universe's,
pippi	pippi,
knyta	tie,
grönland	greenland,
producera	produce,producing,
vattnets	the water's,
fysiologi	physiology,
protoner	protons,
hjärta	heart,
linjerna	routes,lines,
stratton	stratton,
producerad	produced,
modet	the fashion,courage,fashion,
medvetna	aware,conscious,
kommunistisk	communistic,
pennsylvania	pennsylvania,
breda	wide,
hårdvara	hardware,hardwere,
without	without,
nordkoreas	north coreas,
medellivslängd	life expectancy,
lyckan	the happiness,happiness,
helsingfors	helsingfors,helsinki,
listorna	menus,the lists,
kommentarer	comments,
actress	actress,online,
ekologiska	ecological,
enligt	according (to),
allmän	allman,
harrison	harrison,
lyckas	successful,succeed,
leta	check,
utvinns	extracted,
tim	h,
rose	rose,
regent	regent,
rosa	pink,rosa,
utbyte	yield,
utsläpp	emission,emissions,
lett	resulted,
utvinna	extract,
pendeltåg	commuter,
delstat	land,
feminism	feminism,
ross	ross,
riket	kingdom,whole country,
vampyren	the vampire,
delhi	delhi,
virginia	virginia,
uppslagsordet	entry word,lexical entry; word,
kille	guy,
lösas	solved,
inflation	inflation,
vampyrer	vampires,
afrikas	africa's,
kennedy	kennedy,
patrick	patrick,
anföll	attacked,
verksamheten	the work,activity,
madrid	madrid,
teorin	theory,
passera	pass,
latinet	latin,
alkoholer	alcohols,
verksamheter	activity,
försvarare	defenders,defender,
tiders	days',times,time's,
fiktion	fiction,
inspirerades	(was) inspired,inspired,
sitta	sit,
stopp	stop,
härledas	derived,
lärda	scholars,savants,
legat	formed,layed,
uppbyggnad	construction,structure,
storhetstid	heyday,
willy	willy,
football	football,
servrar	servers,
und	und,
geografi	geography,
genom	through,
lyckades	succeeded,
korrekt	proper,
tyska	german,
tyske	german,
förbindelser	connections,relations,
on	on,
om	of,for,
indianska	red indian,amerindian,native american,
spelet	the game,
of	of,
artiklar	items,
stand	stand,
nåddes	reached,
befäl	command,
koppling	clutch,connection,
ansträngningar	effort,
tolkning	interpretation,
burton	burton,
befinna	be,
trådlös	wireless,
fisk	fish,
valley	valley,
serbien	serbia,
förrän	until,
genomfört	carried out,carried through,
flyga	fly,
uppåt	raised,up,
ingredienser	the ingredients,ingredient,
koenigsegg	koenigsegg,
manuskript	manuscript,script,
värre	worse,
taylor	taylor,
felix	felix,
närmast	nearest,
fjorton	fourteen,
tjorven	tjorven,
ökning	increase,
köpenhamn	copenhagen,
många	many,
roses	roses,
mötley	mötley,
regissör	director,
babylon	babylon,
bredare	wider,broad,
separata	separate,
grupp	group,
sällskapet	the company,
symbol	symbol,
erövring	conquest,
missbruk	addiction,abuse,
vinnaren	winner,the winner,
observatörer	observers,
symtomen	the symptoms,
villkor	conditions,condition,
distriktet	district,
calle	calle,
oftast	usually,most often,
erfarenhet	experience,
all	any,
ali	ali,
separat	seperate,
samhället	the society,society,
konsekvent	consistency,
samhällen	societies,
utomliggande	external; ex-territorial,outlying,
sakrament	sacrament,
plikter	duties,
uppdrag	missions,
persiska	persian,
ron	ron,
brottet	offense,
ögonen	eyes,the eyes,
påstående	claim,
program	application,
cykeln	there are two meanings in the context - cycle and bicycle,
kvar	left,
löper	runs,at,
färgerna	colors,
liter	liters,
litet	small,
ansluter	connects,
song	song,
far	father,
fas	phase,
fat	barrel,
runtom	throughout,around,
fan	devil,
sony	sony,
liten	small,
unionens	the union,
tjeckiska	czech,
choklad	chocolate,
helvetet	hell,
list	cunning,
hallucinationer	hallucinations,
förtryck	opression,
lisa	lisa,
iran	iran,
hitta	see,come up, find,
grekland	greece,
ted	ted,
istiden	ice age,the ice age,
tex	e.g.,
design	design,
usama	osama,
enklaste	easiest,
sun	sun,
vaginalt	vaginal,
kinesiska	chinese,
version	version,
sur	acidic,sour,
mördades	was murdered,murder was,
guns	guns,
fäste	bracket,attachment,
christian	christian,
dottern	the daughter,
upptäcka	detection,
regerade	reigned,
avrättades	executed,
leeds	leeds,
fjärdedel	quarter,fourth,
upptäckt	discovered,
norden	scandinavia; (nordic area; region),north,
vilkas	whose,
upptäcks	is discovered,
råder	advises,is,
folktro	folklore,
soloalbum	solo album,
kärnvapen	nuclear,
tillhörde	belonged to,
magnitud	magnitude,
arabemiraten	united arab emirates,uae,the arab emirate,
nyfödda	newborn,
snus	snuff,
uppkomst	origin,onset,
kategorispelare	category player,
filmerna	films,
stöd	support,
syfte	purpose,
smak	taste,
socialdemokraterna	members of the social democracy,social democratic,
anarkism	anarchism,anarchy,
succé	succession,
kommittén	committee,
branden	the fire,
autonom	autonomic,
bekräftade	confirmed,
genomsnittliga	average,
israel	israel,israeli,
permanenta	permanent,
alltid	always,
glas	glass,
hålet	hole,
floyd	floyd,
glad	happy,
östra	eastern,
naturligt	natural,
godkänt	approved,pass,
decenniet	decade,
gatorna	the streets,
decennier	decades,
kryddor	spices,
förhåller	relate,
brown	brown,
bosatt	resident,lived,
huvudort	main town,
elektrisk	electric,
historiskt	historically,
brittisk	british,
satanism	satanism,satanic,
fått	with,
härstamning	lineage,descent,
välgörenhet	charity,
indelade	divided,
rocksångare	rock singers,
taget	time,
böhmen	bohemia,
tagen	taken,
fötterna	the feet,
ångest	anxiety,anguish,
fötts	borned,
atomer	atoms,
regnar	rains,
anarkistiska	anarchistic,
praktiska	practical,
bildade	formed,
tsar	czar,
homosexuella	homosexual,gay,
grande	grande,grand,
greklands	greek gloss,greece's,greek country,
längs	along,
avvisade	rejected,
sträckte	extended,
emmanuel	emmanuel,
mission	mission,
australien	australian,australia,
längd	length,
länge	long,
grupper	groups,
islam	islam,
rike	kingdom,
rika	rich,
rikt	target,rich,
österrikeungern	oster kingdom hungary,
prag	prague,
stephen	stephen,
argentina	argentina,
jämte	together with,
fenomenet	phenomenon,
kategorieuropeiska	european category,europe category,
förebyggande	preventing,preventive,
number	number,
kärna	core,quarks,
postumt	posthumous award,posthumously,
landborgen	the ridge,
marcus	marcus,
försöken	attempts,
forna	former,
slidan	the vagina,vaginal,
journalister	journalists,
försöker	try,
principer	principals,
nervosa	nervosa,
betyg	grades,
hawaii	hawaii,
konstnärlig	artistic,
aldrig	never,
sätt	way,
stenar	stones,blocks,
ollonet	penis head,glans,
därvid	thus; thusly; then,therewith,
väg	way,
kvinna	woman,
väl	selecting,good,
vän	van,
benjamin	benjamin,
poliser	police (-men; -women),
ökad	increase,
islamistiska	islamic,islamist,
beräknades	estimated,
ökat	increased,
spelades	filmed,
ökar	increases,
polisen	police,the police,
faller	fall,
fallet	case,the case,
stavningen	spelling,the spelling,
konsumtionen	the consumtion,consumption,
fallen	cases,
aminosyror	amino acids,
filosofins	philosophy,the philosophy,
heinz	heinz,
colombia	colombia,
pablo	pablo,
bland	inter,
blanc	blanc,
story	story,
infört	introduced,
misslyckas	fail,
stort	large,big,
storm	storm,
brasiliens	brazil's,
ecuador	ecuador,
familjerna	families,
mikael	mikael,
gränser	borders,frontiers,
hotel	hotel,
framtiden	future,
hotet	the threath,the threat,threat,
fattigaste	the poorest,poorest,
två	two,
besökare	visitors,
siffra	number,figure,
king	king,
illegala	irregular,
matcherna	the games,games,
direkt	direct,
mån	concerned,mon,
pjäsen	piece,
dans	dance,
guden	god,the god,
stjärnan	star,
kategorin	the category,
klubb	club,
anläggningar	plants,facilities,
kusin	cousin,
tilldelas	assigned,
tabell	table,
omskärelse	circumcision,
slåss	fight,
divisionen	division,
wilson	wilson,
dialekt	dialect,
jämförelsevis	comparative,
judas	judas,
unge	young,
folkgrupper	ethnic groups,
electric	electric,
dagliga	daily,
naturvetenskapliga	scientific,
dagligt	daily,
industrialiserade	industrialized,
europarådet	european council,
sånger	songs,
mineral	mineral,
windows	windows,
salt	salt,
influensan	the influenza,flu,
statsskick	government,
kosovo	kosovo,
tjugo	twenty,
ursprungliga	original,
kolonialism	colonialism,
tilly	tilly,
månen	the moon,man,
förening	union,
beräkningar	calculations,
canaria	canaria,
grace	grace,
moses	moses,
hit	here,
hiv	hiv,
stormakterna	great powers,
vardera	either,each,
b	b,
jobbade	worked,
händer	happens,
himmler	himmler,
utvidgade	expanded,
mediciner	medicines,
avtal	agreement; deal,
tidszon	time zone,
vincent	vincent,
norrköping	norrköping,
poäng	score,point,
utsatt	exposed,
bars	bar,
etiopien	ethiopia,ethiopian,
art	kind,art,
bart	bart,
arv	heritage,
butiker	stores,
bara	only,
are	are,
förtroende	trust,
flyttade	moved,
stjäla	steal,stealing,
arm	arm,
barn	child,
bortsett	except,
planeras	planned,
planerar	is planning,plan,planned,
inga	not,
invaldes	was elected,
planerad	planned,
oerhörd	tremendous,
verksamhet	activity,
intäkter	revenues,incomes,
uppkom	arose,
godkändes	approved,
vätet	hydrogen,the hydrogen,
tiderna	the times,
startades	started,
roman	novel,
klassificeras	classified,
hypotesen	the hypothesis,
lära	lara,get to know,
smith	smith,
vidare	further,furthermore,
stärktes	strengthened,
belägna	located,disposed,
besegrade	defeated,
östtyskland	east germany,
utifrån	from,
hypoteser	hypotheses,hypothesis,
ps	ps,p.s,p.s.,
java	java,
göteborg	gothenburg,
personalen	personnel,the staff,
kungafamiljen	the royal family,
pc	pc,personal computer,
byxor	pants,
ska	will,
ph	ph,
pi	pi,
flight	flights,flight,
togs	taken,
publiken	audience,
sydafrikas	south africa's,
rättigheterna	rights,
gården	courtyard; house; farm (-house),
konflikter	conflict,
konflikten	the conflict,conflict,
sådan	such,kind of,
inspelningar	recordings,
generationer	generation,
ris	rice,
rik	rish,rich,
skeppen	the ships,
demografi	demography,
tidpunkten	the time,
ideologier	ideologies,
sjunkit	decreased,
förföljelse	persecution,
torbjörn	torbjörn,
spears	spears,
låtit	had,ordered,
skeppet	the ship,
byar	villages,
skåne	skåne,
berömd	famous,
experimenterade	experimented,
berömt	famous,
vinklar	angle,angles,
finansiera	fund,
italiensk	italian,
sjunga	sing,
edge	edge,
kyrkans	the church's,
alfabet	alphabets,
uttalande	statement,
kontinentala	continental,
komplett	complete,
konstitution	constitution,
påverkade	influenced,affected,
remmer	remmer,
namnet	name,the name,
folkräkning	head count,public shaving,
minoriteter	minorities,
bostad	property,
omedelbar	instant,
försvunnit	disappeared,
skall	is,
centralasien	central asia,
idé	regard,
emigrerade	emigrated,
skala	scale,
rastafarianerna	the rastafarian,
begravdes	buried,
användas	used,
stoppade	stop,
upplevelse	experience,
exakt	precise,accurately,
våldsamma	violent,
banbrytande	groundbreaking,
sammansättning	composition,
hittades	was found,
hittas	found,
hittat	found,
minskning	reduction,decrease,
norrut	north,
sjöfart	sea voyage,maritime,
kongo	congo,kongo,
global	global,
flottan	navy,
thailand	thailand,
låtarna	the songs,
ungefär	approx.; approximately,
höjden	height,
grekerna	greeks,
statyn	the statue,
frälsning	salvation,
fungera	act,
anne	anne,
anna	anna,
höjder	heights,
turism	tourism,
diamant	diamond,
palmes	palme's,
ställningen	position,
tävlade	competed,
lånat	borrowed,
anklagades	accused,
bayern	bavaria,bayern,
judendom	judaism,
kostnaderna	costs,the costs,
grundläggande	because lag of,fundamental,
påtryckningar	pressure,
tätt	tight,tightly,
vägarna	paths,roads (roadways),
täta	close,
socialistisk	socialistic,
oktoberrevolutionen	the october revolution,
genomföras	carried out,be performed,carry out,
reglerna	rules,rules; regulations,
hållet	attached via,cohesive,
inblandade	involved,
km²	km2,
håller	halls,
uppvisar	shows,
long	longitude,long,
bruk	use,
laila	laila,
ateister	steister,
delning	division,pitch,
rasade	collapsed,
regionen	the region,region,
sköter	handles,handle,
kritikerna	critiques,
delta	participate,delta,
tidigast	the earliest,
junior	junior,
medeltidens	medieval,
anklagelser	allegations,
planeternas	the planets',
angels	angels,
styrande	rulers,
variant	variant,
utrikespolitik	forgein policy,
erövrades	(was) conquered,
guyana	guyana (name),guyana,
tolka	interpret,
fick	got,was,
z	z,
svenskspråkiga	swedish-speaking,
ägdes	owned,
singlarna	the singles,simglama,
tidpunkt	time,
däribland	among them,including,
graham	graham,
veckorna	weeks,
rainbow	rainbow,
stadion	stadium,the stadium,
möten	moten,
liechtenstein	liechtenstein,
psykoterapi	psychotherapy,
högst	maximum,
hanen	the cock,male,
urval	selection,
skyddas	skyas,
skyddar	protects,
sutra	sutra,
beräknar	calculates the,computes,
tittarna	viewers,
medina	medina,
konvertera	conversion,
jugoslaviska	jugoslavian,
modernismen	modernism,
oväntat	unexpectedly,
underlättar	facilitates,
vice	vice,
europeiska	european,
målvakten	the goalkeeper,
microsoft	microsoft,
nasa	nasa,
karma	karma,
lagstiftning	regulation,
europeiskt	european,
nash	' nash,
förhandla	negotiate,
psykologi	psychology,
beträffande	on,
kanal	channel,
steve	steve,
jimi	jimi,
låter	let,
moseboken	genesis,
norrköpings	norrköpings,
simon	simon,
fortfarande	still,
generella	overall,general,
hinduism	hinduism,
fotnoter	footnotes,
varierar	vary,
vapen	weapons,
kategoritvseriestarter	category television series starts,
varierat	varied,
kommitté	committee,
tvinga	force,
historikern	the historian,
demokratiskt	democratic,
äta	eat,
byggt	built,
noter	notes,
öron	anxiety,ears,
julius	julius,
utanför	outside,
melodier	melodies,
byggd	built,
bygga	building,
indirekt	indirect,
skadad	damaged,
åtta	eight,
århundradet	century,
skadan	the hit,the damage,
influerad	influenced,
skadas	damaged,
västlig	western,
konstant	constant,
folk	public,
dramatiskt	dramatically,
assisterande	assisting,
kris	crisis,
judy	judy,
krig	war,
dramatiska	dramatic,
koloni	colony,
hdmi	hdmi,
producenten	the producer,producer,
turismen	tourism,the tourism,
producenter	producers,
diamanter	diamonds,
åtgärder	measures,
expansion	expansion,
astrid	astrid,
fauna	fauna,
ukraina	ukraine,
metro	metro,
innehar	holds,
innehav	possession,
springsteens	springsteens,
plattan	plate,the plate,
fortsätter	continues,continue,
populärkulturen	popular culture,
tjänar	earns,
zlatan	zlatan,
reda	find out,out,find our,
gemenskap	fellowship,community,
redo	ready,prepared,
varpå	thereafter,
from	from,
bestämmelser	conditions,
usa	the usa,
fel	faults,
sevärdheter	attractions,
vikingar	vikings,
upplöstes	dissolved,
källorna	source,the sources,
inlandet	inland,
öppnat	opened,opening,
andliga	spiritual,
penis	penis,
införande	introduction,
hindrade	preventing,prevented,
vägrade	refused,
fungerar	functions,works,
reguljära	regular,
beskriva	describe,
automatiskt	automatic,
beskrivs	described,
tas	is,is taken,
platser	points,
crick	crick,
platsen	the place,site,
tag	while,
hilton	hilton,
tal	speech,
kanadensiska	canadian,
sir	sir,
beyoncé	beyonce,beyoncé,beyoncè,
six	six,
brian	brian,
sig	to,
undantaget	except,
sin	its,
väpnad	armed,
kontroversiellt	controversial,
förekommande	occuring,where,
oavsett	whether,regardless; whether; irrespective of,
tack	thanks,
religiös	religious,
lätta	lighten,
kontroversiella	controversial,
eritrea	eritrea,
light	light,
centralorter	centers,
framförts	forward,
företag	company,companies,business,
jolie	jolie,jolies,
besegrat	defeated,
mekka	mecca,mecka,
blandad	blended,
skapande	building,creative,
företrädare	representatives,
förklaras	explained,
elit	elite,
blandat	mixed,
karlstad	karlstad,phoenix,
blandas	mixed,
spotify	spotify,
listan	the list,
uppmärksammad	attention,
terriers	terriers,
befolkning	population,
byn	village,
återvänt	atervant,returned,
försvar	defence,defense,
datorn	the computer,pc,
uppmärksammat	attention,noticed,
carola	carola,
cypern	cyprus,
betalade	paid,
underjordiska	underground,
omedelbart	immediately,immediate,
östtimor	east timor,
redovisas	shown,
satelliter	satellite,
exempelvis	e.g.,
växande	growing,
konungariket	kingdom,
vidta	take,
studios	studios,the studio's,
australiska	australian,
barnets	the child's,
byter	changing,changes,
kvarteret	quarter,the neighborhood,
säsongen	season,
arterna	species,
kritik	critisism,critique; criticism,
förbjuda	forbid,ban,
uggla	owl,
minskad	reduced,
hantverkare	craftsman,
fiktiva	fictitious,romantic,
svar	answer,response,
bål	prom,torso,
nobelpristagare	nobel laureate (-s); nobel prize winner (-s),
minskat	has decreased,
centralamerika	central america,
minskar	decrease,diminishing,
förutsättningar	prerequisites,(pre-)conditions,condition,
hörs	heard,
ifrån	off,
hjälpt	helped,
vulkanutbrott	vulcano eruption,
utmärker	characterizes,characterized,
höra	hear,know,
hjälpa	helping,
studioalbumet	studio album,
philip	philip,
domare	judge,
hörn	corner,
fotbollslandslag	football team,national football team,
gångna	past,
anslutning	connection,
tyst	quiet,silent,
kortare	shorter,
g	(g),
barns	childrens,
adrian	adrian,
tysk	german,
rudolf	rudolph,
belagt	coated,
revolutionens	revolution,the revolutions,
isbn	isbn,
värsta	worst,
regenter	monarchs,
skyddade	protected,
nätverk	network,
enkelt	easy,
åtskilliga	several,
fågelhundar	bird dogs,
meddelanden	messages,
omfattning	extent,
misslyckande	failure,
sankta	sankta,
diskutera	discussed,
rösträtt	vote,right to vote,
valde	selected,chose,
valda	chosen,
vingar	wings,
juli	july,
vind	wind,
dödligheten	mortality,
bevarade	preserved,
franska	french,
holland	holland,
franske	the french,french,
birgitta	birgitta,
franskt	french,
tyskarna	the german,
farliga	dangerous,
romarna	the roman,the romans,
cohen	cohen,
flyttar	move,
avgörs	determined,
blir	become,is,
farligt	dangerous,
ringen	ring,
intervju	interview,
storbritannien	great britain,uk,
byggas	prevented,build,
uppfann	invented,
lopp	course, passage,
kristi	kristi,christ,
betydligt	significant,
centra	center,
centre	centre,
intogs	was taken,was captured,
väntat	expected,
staternas	the state's,
öken	ok,desert,
förbundsrepubliken	the federal republic,federal republic of,
regeringschef	head of government,government,
miljontals	millions,
enbart	only,
generna	genes,the genes,
kategoriamerikanska	u.s. category,
movie	movie,
moberg	moberg,
uefa	uefa,
blandade	mixed,
funktionella	functional,
debatt	debate,
julafton	chistmas eve,
pastoral	pastoral,
angående	reference,
filmen	film,
rösten	voice,rust,
filmer	movies,
röster	votes,
piano	piano,
allmänhet	in general,public,
träffa	see,
gränsar	adjacent,
heta	hot,be named; be called,be called,
gudar	gods,
linje	line,
närstående	relatives,kindred,
samtycke	consent,
städer	urban,
begäran	request,
torka	dry,
mestadels	most of the time,mostly,
kvinnorna	the women,
nationernas	the nations,
rikare	richer,
motståndare	opponents,opponent,
theta	theta,
funktion	function,
upplysning	the enlightenment,enlightenment,
praktisk	practical,
sydstaterna	southern states,southern united states,
swift	swift,
jon	jon,
sångaren	singer,the singer,
styrdes	ruled,
allsvenskan	headlines,allsvenskan,
påtagligt	considerably,markedly,
utvecklingen	the development,
teoretiker	say,theorists,
kolhydrater	carbons,carbohydrates,
april	april,
västerländsk	western,
republikens	republic's,republic,
bronx	bronx,
förespråkare	spokesman,proponent,
betecknar	represent,
betecknas	labelled,
exakta	exact,
korruption	corruption,
wall	wall,
publicerad	published,
walt	walt,
cirka	about,
utsedd	appointed,
innebära	mean,
publiceras	will be published,
framträdanden	appearances,
publicerat	published,
klara	clear,
hindu	hindu,
bbc	bbc,
beskrivning	description,
månar	moons,
klart	finished,done,
strindbergs	strindberg's,strindberg,
ständig	constant,
naturtillgångar	natural resources,
mike	micke,mike,
liverpool	liverpool,
nickel	nickel,
klassen	klasses,
turneringen	the tournament,
dominera	dominate,
lutherska	lutheran,
försvann	disappeared,
hms	hms,
fortsättningen	remain,the continuation,
neutrala	neutral,
deklarerade	declared,
antogs	adoption,was assumed,
godkännande	approval,
bråk	brawl; fight,fraction,
officiell	official,
största	biggest,
anpassa	adapt,
will	will,
fördelade	divided,
wild	wild,
madeleine	madeleine,
kommande	upcoming,
explosionen	the explosion,
uppfattning	view,
gemensamt	single,in common,
själ	soul,
syftar	refers,refer,
motiv	subjects,
röra	move,
uppstå	develop,occur,
halv	half,
buddhism	buddhism,
pojkar	boys,
samband	connection,
inch	inches,
skickade	sent,
gett	gave,
kustlinje	coastline,
mottagande	host,
övervägande	the predominant,
romeo	romeo,
romer	roma,
student	student,
raka	straight,
rätt	steering wheel,
misstag	error,
klubbar	clubs,
vilar	rests,
banden	bands,
undersökningar	studies,studies',
närma	approach,move closer,approximate,
ekosystem	ecosystem,eco system,
övertyga	convince,
bandet	band,
organisationens	organization,
hårdrocken	hard rock,
lön	salary,wage; salary,
biologisk	biological,
singeln	single,singeln,
mfl	etc,etc.,
möjligheter	potential,
uppkommer	arises,arises; generated,
rachels	rachel's,
erfarenheter	experiences,experience,
högskolor	colleges,
patrik	patrik,
miljöer	environment,environments,
antisemitism	antisemitism,
rocken	the rock,rock,
brutit	cut; break,
mytologiska	mythological,
jarl	earl,
alldeles	completely,altogether,
hoppa	skip,
sky	sky,
rättsliga	justice,
engelsk	english,
ske	be,
resultat	result,
fyller	turns,turn; fill,
sanskrit	sanskrit,
psykoser	psychoses,psychosis,
älska	love,
know	know,
press	press,
psykosen	psychosis,
säljs	sold,
georges	georges,
miami	miami,
djupa	deep,
huruvida	whether,
sälja	sell,
gorbatjov	gorbachev,
globalt	globally,global,
finansieras	financed,funded,
djupt	deep,
säkra	safe,
juni	june,
tjeckoslovakien	czechoslovakia,
handeln	trade; commerce,
efterfrågan	demand,
aktier	share,stock,
handels	commercial,trade,
försvinna	disappear,
empire	empire,
skandinavien	scandinavia,
använts	used,
planering	planning,
trianglar	with triangles,
gammalt	old,
risker	risker,
setts	observed,
personligen	personally,
stieg	stieg,
låten	the song,song,
sjunker	flag,sinks,
markera	mark,
utsöndras	secreted,
uppvärmning	heating,
mitt	my,
slut	end,
dateras	dates,
sommarspelen	summer games,summer olympics,
ljung	heather,
låna	borrow,lana,
koalition	coalition,
substantiv	noun,
tillräcklig	sufficient,
bestämma	determining,
oberoende	independent,
avsnittet	section,episode,
saken	the thing,the matter,
saker	items,
reaktionerna	the reactions,reactions,
mäta	feeding,
främre	forward,
egna	own,
floder	rivers,
stanna	stop,
avrättade	executed,
tillbringade	spent,
mäts	is measured,
en	a,
floden	the river,
mätt	dull,
flyger	flies,flying,
stressorer	stressors,
glukos	glucose,
folkpartiet	peoples party,liberal party,
konstruktion	structure,
van	van,
flamländska	flemish,
upprättas	established,
vad	as,what,
smeknamnet	nickname,
mäter	measure,
var	was,
regisserad	directed,
vacker	beautiful,
nordamerikanska	north american,
granne	neighbour,
hundratal	100,hundred,
ingått	been part of,entered,entered into,
krigsslutet	end of the war,
stadens	the citys,city's,
karta	map,
rybak	rybak,
tema	theme,
missnöjet	discontent,
jenny	jenny,
problemet	the problem,
stormakter	world powers,
eu	eu,
runor	runes,
resultera	result,
året	the year,all year,
illinois	illinois,
ursprunget	origin,the origin,
åren	the years,years,
serbiska	serbian,
tolkas	interpretation,
tolkar	interprets,
shakespeares	shakespeare's,shakespeare,
tvfilm	tv-movie,
mankell	mankell,
ställningar	standings,notions,
margaret	margaret,
markant	considerably,markedly,
nödvändigtvis	by necessity,
knappast	hardly,dead,
bysantinska	byzantine,
simpson	simpson,
tidning	journal,
