vanligast	most usual,most common,
nordisk	nordic,
uppemot	almost,
stammarna	tribes,
arternas	the species,
elva	eleven,
invandrare	immigrant,
hållas	be held,
slå	hit,
albumen	the albums,
hermann	hermann,
vann	won,
lyckats	succeeded,
dela	divide,
syrgas	oxygen,
upptar	occupies,
skicklig	skillful,
statlig	government,
medelhavet	mediterranean sea,
haber	haber,
befogenheter	authorities,
urskilja	discern,
sture	sture,
sammansatta	composed,
ungerns	hungrarys,
hanar	males,
upprätthåller	maintains,maintaining,
åsikten	the opinion,
punkt	point,
österrike	austria,
hårda	hard,
biografi	biography,
vägrar	refuses,refuse,
filosofen	the philosopher,
motståndsrörelsen	the resistance,
regnskog	rain forest,
analytisk	analytical,
bipolär	bipolar,
kids	kids,
demokratier	democracies,
naturen	the nature,
blåser	blowing,
miljarder	billions,
karin	karin,
systematiska	systematical,
biskop	bishop,
välkänd	well known,
systematiskt	systematic,
ansluta	connect,
dna	dna,
strikt	strict,
fuktiga	damply,
 mm	millimeter,
dns	dns,
fuktigt	moist,
musik	music,
befolkningstillväxten	the population growth,the growth of population,
mercurys	mercury's,mercurys,
holm	holm,
politiker	politician,
bulgariska	bulgarian,
teman	themes,
ofta	often,
vännen	the friend,
befolkningsutveckling	population development,
vågen	the wave,
stommen	the foundation,
passagerare	passenger,
kapitalismen	capitalism,
hon	she,
kallare	colder,
pågick	lasted,
typen	the type,type,
fylla	fill,
inrikes	domestic,
barbro	barbro,
sedd	seen,
turkiet	turkey,
sankt	sankt,
typer	types,
hisingen	hisingen,
grekiska	greek,
hemsida	homepage,
hemlandet	the home country,the homeland,
wind	wind,
vart	each,
varv	dockyard,
ormar	snakes,
dalí	dali,
organismen	the organism,
varg	wolf,
vara	be,
mabel	mabel,
varm	warm,
publicerade	published,
målade	painted,
assyriska	assyrian,
fil	master of,
avgå	resign,
myntade	coined,
hänga	hang,
närliggande	nearby,
silver	silver,
utvecklat	evolved,
utvecklar	develops,
vattenånga	steam,
terrorister	terrorists,
debut	debut,
utveckling	development,
tillgängligt	available,
utvecklad	developed,
tillgängliga	available,
angola	angola,
serier	comics,
allan	allan,
kontroverser	controversies,
serien	the series,
truman	truman,
varken	either,
george	george,
försökt	tried,
förändringar	changes,
debatter	debates,
anarkister	anarchists,
underordnade	subordinates,
sannolikt	probable,
att	that,
sysselsätter	employs,
malmös	malmö's,
givetvis	naturally,
grannlandet	the neighbouring country,
östberg	Östberg,
tecknade	drew,
förespråkar	advocate,
xis	the eleventh's,
master	master,
ära	glory,
bitter	bitter,
bokstäverna	the letters,
förmögenhet	wealth,
placerade	placed,
nirvana	nirvana,
påverkad	influenced,affected,
ahmed	ahmed,
skatter	taxes,
upphov	origin,source,
stormaktstiden	great power period,
påverkan	impact,influence,
tree	tree,
gator	streets,
nations	nations,
trey	trey,
varje	each,
utformningen	the layout,
tretton	thirteen,
obligatorisk	mandatory,
försörja	support,
assistent	assistant,
kriterierna	criteria,
boston	boston,
filosofisk	philosophic,
joakim	joakim,
trakten	the region,region,
normalt	normally,
östeuropa	east europe,
skaffa	obtain,
förhärskande	prevailing,
hjälpmedel	aid,
bedrivs	conducted,
konserthus	concert hall,
gallagher	gallagher,
anteckningar	notes,
bedriva	prosecute,
thriller	thriller,
övertog	overtook,
singer	singer,
arkitektur	architecture,
hämnd	revenge,
camp	camp,
utmärkande	distinguishing,
förlorar	loses,
förlorat	lost,
grovt	heavy,
passerade	passed,
singel	single,
tänkte	thought,
majs	corn,
anorektiker	anorectic,
konkret	concrete,
legitimitet	legitimacy,
teater	theater,
buss	bus,
övergår	surpasses,
sekulär	secular,
bush	bush,
lastbilar	truck,
tillståndet	the state,
årsdag	anniversary,
upprätta	establish,
metoden	the method,
dansk	danish,
plats	place,
bensin	gasoline,
innebörd	meaning,
spänning	voltage,
kallt	cold,
sköta	operate,
utgåvan	the edition,
uppgift	task,
genomsnittet	average,
statschef	head of state,
kalla	cold,
blev	became,
etik	ethics,
flagga	flag,
skulle	would,
skriva	write,
arlanda	arlanda,
best	best,
hedersdoktor	honorary degree,
manson	manson,
wikipedia	wikipedia,
sista	last,
ringa	call,
rollen	the role,
lanserades	was launched,
tilldelades	awarded,
kommunikation	communication,
världsturné	world tour,
roller	roles,
tillämpar	practice,administers,
tillämpas	applied,
pitt	pitt,
anordnas	arranged,
nordiskt	nordic,
genus	genus,
logik	logic,
summan	the sum,
igelkotten	the hedgehog,
armén	the army,
herr	mister,
ana	feel,
avgörande	settling,
fri	free,
tiotusentals	tens of thousands,
operationer	operations,
socialistiskt	socialistic,
årtionde	decade,
stadium	stage,
arbetslösheten	unemployment,
verktyg	tools,
barndom	childhood,
life	life,
café	café,
ändrade	changed,
arkiv	archive,
närvarande	present,
dave	dave,
kometer	comets,
chile	chile,
övergripande	general,
chili	chili,
parterna	parties,
intag	intake,
uttryck	expression,
frankrikes	frances,
castro	castro,
organisera	organize,
kontraktet	the contract,
tintin	tintin,
brister	inabilities,
förföljelser	pursuits,persecutions,
desto	ever,
player	player,
tänkare	thinker,
bristen	lack of,
slag	kinds,
madonna	madonna,
tät	compact,sealed,
serbisk	serbian,
tillhandahåller	provides,
vrida	twist,
foton	photos,
funktionen	the function,
josef	josef,
topp	top,
emi	emi,
föras	be brought,
synder	sins,
tung	heavy,
zeeland	zeeland,
kampanj	campaign,
gudinnan	the godess,
grundlag	constitution,
försvarade	defended,
snö	snow,
köra	drive,
capitol	capitol,
dödsoffer	casualty,death victim,
norsk	norwegian,
körs	driven,being driven,
utrotning	extinction,
kommunal	communal,municipal,
döda	dead,
matteus	matteus,
vetenskapsmän	scientist,
bnp	gdp,
uppgörelse	agreement,
hette	named,
lunginflammation	pneumonia,
hav	seas,ocean,
underliggande	underlying,
svensson	svensson,
livsstil	lifestyle,
dagar	days,
uppmärksammade	observed,
county	county,
bobby	bobby,
alice	alice,
kust	coast,
residensstad	city of residence,county seat,
sebastian	sebastian,
ola	ola,
företräder	representing,
people	people,
parlamentarisk	parliamentary,
delade	split,
kulmen	the acme,
fot	foot,
varierande	varied,varying,
utses	is appointed,
akademi	academy,
idéer	ideas,
myndigheter	authorities,
annan	another,
stefan	stefan,
påminner	reminds,
hörde	heard,
olympiska	olympic,
möjligheterna	the possibilities,
myndigheten	the authority,
annat	other,
nixon	nixon,
hänt	happened,
delvis	partially,
psykiska	mental,
marshall	marshall,
som	as,which,
sol	sun,
lagliga	legal,
psykiskt	psychic,
nova	nova,
säkerhetspolitik	safety policy,
 miljoner	millions,
offer	victim,
öppen	open,
förhållanden	relationships,
öppet	open,
verde	verde,
tigern	the tiger,
avsevärt	substantially,
drabbat	affected,
gymnasiet	high school,
drabbar	affect,troubles,
polska	polish,
syften	purpose,
pest	plague,
moderna	modern,
föregångare	predecessor,
konung	king,
lunds	lund's,
låtar	songs,
krävde	demanded,
ericsson	ericsson,
dotter	daughter,
protester	protests,
republik	republic,
olja	oil,
reggae	reggae,
avskaffades	was abolished,
bostadsområden	residential areas,
jamaicanska	jamaican,
blått	blue,
vintrarna	the winters,
modell	model,
transporter	transports,
tävling	competition,
sällan	rare,
förtjust	delighted,
trettio	thirty,
time	time,
skatt	tax,
erkände	acknowledged,
ost	cheese,
uppgifter	tasks,data,
stödjer	supports,
uppgiften	the task,
atombomben	the nuclear bomb,
traditionell	traditional,
inkomst	income,
machu	machu,
vet	know,
fängelset	prison,
intresserade	interested,
grön	green,
vem	who,
bosnien	bosnia,
musikstilar	music genres,
choice	choice,
individen	the individual,
skillnaderna	the differences,
kompositörer	compositors,
inhemska	native,
saab	saab,
jämnt	even,evenly,
jämna	even,
firandet	the celebration,
jämföras	compared,
köp	purchase,
kunskapen	the knowledge,
axel	axel,
kön	gender,sex,
kunskaper	knowledge,
provinserna	the provinces,
galileo	galileo,
vintertid	winter-time,
katten	the cat,
huvudsakliga	main,
studien	the study,
genomgående	consistently,
bärande	leading,
studiet	the study,
studier	studies,
santa	santa,
sprids	spreads,
samlat	gathered,
positiva	positive,
änglar	angels,
sprida	spread,
positivt	positive,
ställt	taken,put,
dagars	days,
relationerna	the relationships,
ställe	place,
ställa	set,
grönt	green,
gröna	green,
påvisa	show,
stigande	rising,
missförstånd	misunderstanding,
locke	locke,
släktskap	kinship,
inkluderade	included,
kretsar	circles,
korta	short,
milda	mild,
årligen	annually,
begick	commited,
svenskan	swedish,
européer	europeans,
riksdagen	the parliament,
gigantiska	gigantic,
kungens	the king's,
löpande	running,
svart	black,
nyligen	recently,
data	data,
epost	email,
portugisiska	portuguese,
bergarter	rock types,rocks,
undervisning	education,
ss	ss,
st	saint,
sk	so called,
sm	swedish championship,
sa	said,
vika	fold,
se	see,
resulterar	result,
vintrar	winters,
resulterat	resulted in,
kong	kong,
antingen	either,
allvarligt	serious,
ersätta	replace,
ingvar	ingvar,
dialekter	dialects,
utsätts	exposed,
jim	jim,
tilldelats	awarded,
turnera	tour,
faderns	the father's,
monopol	monopoly,
personlig	personal,
hos	with,
öppnades	were opened,was opened,
musiken	the music,
matcher	matches,games,
sorter	kinds,
matchen	the game,
kantoner	cantons,
förväxlas	confused,
omöjligt	impossible,
skivkontrakt	record contract,
dominerar	dominates,
runstenar	runestones,
dominerat	dominated,
födelsedag	birthday,
dynamiska	dynamic,
står	standing,
krav	requirement,
kött	meat,
riktigt	real,
bly	led,
sjuka	sick,
densitet	density,
bli	become,
bränder	fires,
internet	internet,
roterar	rotates,
sfären	sphere,
vård	healthcare,
våra	our,
bytt	traded,
byts	replaced,
sålda	sold,
kolonier	colonies,
byta	change,trade,
pund	pound,
punk	punk rock,
artisten	the artist,
gordon	gordon,
gård	farm,
hård	hard,
tsunamier	tsunamis,
hårt	hard,
open	open,
ont	bad,
city	city,
teologi	teology,theology,
råolja	crude oil,
intill	beside,adjacent to,
sjö	lake,
nästa	next,
williams	williams,
vilka	who,
tillräckligt	sufficient,
irakiska	iraqi,
tillräckliga	insufficient,sufficient,
svenskarna	the swedes,
provins	province,
dygn	day,
fiskar	fishes,
kamprad	kamprad,
motståndarna	the opponents,
tankar	thoughts,
sak	thing,
konsekvenser	consequences,
församlingar	parishs,
känslan	the feeling,
allen	allen,
staden	the city,
priserna	the prices,
övriga	others,
takt	rate,
zon	zone,
jefferson	jefferson,
harald	harald,
övrigt	other,
förändringen	the change,
muslimer	muslims,
finlands	finlands,
sekreterare	secretary,
mynt	coin,
religionen	the religion,
forskningen	the science,
driva	operate,
phil	phil,
inledningen	the introduction,
ursprung	root,
rykte	reputation,
kvicksilver	mercury,
drivs	driven,
engagemang	commitment,
olagligt	illegal,
axl	axl,
beckham	beckham,
dimensioner	dimensions,
sjöss	sea,
antalet	number,the number,
stärkte	strengthened,
västsahara	western sahara,
hockey	ice hockey,
belgien	belgium,
inlägg	post,
platta	flat,
undersöka	research,
rörande	concerning,
ländernas	the countries,
artist	artist,
råd	council,
antogs	was assumed,
erbjöds	offered,
vision	vision,
brännvin	schnaps,
snabbare	faster,
behovet	the need,
nederbörden	the precipitation,
skärgård	archipelago,
talman	spokesperson,
ordspråk	proverb,
enhetlig	uniform,
utgörs	consists of,
källa	source,
kritiserade	critisized,criticized,
begränsningar	limitations,
upplever	experience,
utgöra	compose,make up,
kilometer	kilometer,kilometers,
små	small,
anledningarna	the reasons,
screen	screen,
amerikanske	american,
awards	awards,
amerikanska	american,
mariette	mariette,
basisten	basist,the basist,
mans	man's,
rekord	record,
mani	mania,
tillsätts	appoints,
långsammare	slower,
upproret	the upprising,
klimat	climate,
hamnade	landed,
drogs	was pulled,
farfar	paternal grandfather,
bolag	company,
luft	air,
cupen	the cup,
lidit	suffered,
lånat	borrowed,
formen	the form,
formel	formula,
arabiska	arabian,
tillåtet	allowed,
samling	collection,
förstnämnda	first named,
situation	situation,
aston	aston,
bror	brother,
bron	the bridge,
slovenska	slovenian,
nation	nation,
tillåtelse	permission,
blad	leaves,
beteckna	denote,
världsbanken	world bank,
försäkra	make sure,
träffat	met,
ärftliga	genetic,
träffar	meets,
oceanen	the ocean,
ekologi	ecology,
nationalparker	national parks,
brändes	burned,
singapore	singapore,
sägas	is said,
lindgrens	lindgrens,
harris	harris,
senator	senator,
dsmiv	dsm-iv,
händelsehorisonten	the event horizon,
avser	regard,
avses	regard,
summer	sommar,
förluster	losses,
bokförlaget	bokförlaget,
berättelse	story,
koncentration	concentration,
spårvagnar	trams,
höglandet	the highland,
resa	travel,
libyen	libya,
förlusten	loss,
helige	holy,
isen	the ice,
instrument	intrument,
körberg	körberg,
infördes	introduced,
unikt	unique,
regim	regime,
unesco	unesco,
skadade	wounded,
stammar	stutters,
statsreligion	state religion,
tsunami	tsunami,
intet	nothing,
jobbar	work,
nämnas	mentioned,
ursprungsbefolkning	native population,
kännedom	knowledge,
strindberg	strindberg,
institutionerna	institutions,
än	yet,
exil	exile,
katolsk	catholic,
jacksons	jackson's,jacksons,
medlemsstater	member-state,
organisationen	the organization,
herrlandslag	men's national team,
vissa	some,
populationen	the population,population,
digerdöden	the black death,
populationer	populations,
sättas	turn,
förbundskapten	manager,
visst	certain,
ägnar	spend time,spends time,
berger	berger,
upplevelser	experiences,
ronden	round,
berget	the mountain,
nationalencyklopedin	the national encyclopedia,
tillägg	addition,
partiet	the party,
partier	parties,
het	up to date,
förintelsen	the genocide,
philadelphia	philadelphia,
evangeliska	evangelical,
hamnen	the harbour,
hänvisning	reference,
alltså	therefore,really,
bevarat	preserve,
bevaras	are protected,
språkliga	linguistic,
bevarad	kept,
rush	rush,
jamaicas	jamaicas,
kvartsfinalen	quarter finals,quarterfinals,
vinkeln	the angle,
afrodite	afrodite,
förbundsstat	federal state,
age	age,
regimer	regimes,
ac	ac,
redovisas	accounted for,
gustafs	gustafs,gustaf's,
al	alder,
bronsåldern	the bronze age,
beordrade	ordered,
av	of,
håll	ways,
väsentligt	relevant,
federala	federal,
rökning	smoking,
innehåll	content,
svårt	difficult,
belönades	awarded,
avslöjade	revealed,
värt	worth,
koppar	copper,
gifte	married,
kvarstod	remained,
medverkat	participated,
medverkar	contributes,contribute,
forntida	prehistoric,
vinner	wins,
beteckning	label,
decennierna	decades,
original	original,orignal,
renässans	renaissance,
släppt	released,
resor	travels,
elektron	electron,
halsen	the throat,
kammare	chamber,
släppa	release,
likartade	similiar,
norr	north,
skogarna	the forests,
pojkvän	boyfriend,
ullevi	ullevi,
tv	tv,
nederbörd	rainfall,
mildare	milder,
nord	north,
te	tea,
strand	beach,
utländsk	foregin,
sant	true,
djurarter	animal species,species,
borrelia	borreliosis,
muslimska	muslim,
utsåg	declared,
siffrorna	numbers,
smala	narrow,
harry	harry,
språkbruk	parlance,
döttrar	daughters,
påståenden	claims,assertions,
synd	sin,
dödsstraff	death penalty,
utökade	expanded,
skede	period,
givaren	the giver,
övergav	abandoned,
delen	part,
islams	islams,islam's,
hänsyn	consideration,
full	full,
gruppen	the group,
arkeologiska	archaeological,
november	november,
legend	legend,
motstånd	resistance,opposition,
traditionella	traditional,
exklusiv	exclusive,
traditionellt	traditional,
social	social,
oftare	more often,
varelser	creatures,
sena	late,
kommunistpartiet	the communist party,
vid	by,
ordinarie	regular,
vin	wine,
juridiskt	judicial,
kuiperbältet	the kuiper belt,
vit	white,
främja	further,
skapa	create,
biskopen	the bishop,
petroleum	petroleum,
pearl	pearl,
sitter	serve,sit,
dödligt	lethal,deadly,
mora	mora,
fyrtio	forty,
berättade	told,
uppskattas	is appreciated,
uppskattar	estimates,
schweiz	switzerland,
undergång	doom,
inträffade	happened,
medelklassen	middle class,
science	science,
beskyddare	protector,patron,
cykel	bicycle,
kapitalism	capitalism,
läkaren	the doctor,
samväldet	the commonwealth,
nobelpriset	the nobel prize,
säljas	is sold,
nordvästra	northwest,north western,
skadliga	harmful,
mellersta	middle,the middle,
stater	states,
spansk	spanish,
järnvägsnätet	railroad network,
information	information,
vägnätet	road network,
hugo	hugo,
uppfattade	perceived,
ansetts	regarded,
lejon	lion,
riksdagens	the parliament's,the parliaments,
fortsättning	continuation,
kedjan	the chain,
soundtrack	soundtrack,
lanka	lanka,
anklagade	accused,
komplexa	complex,
hållit	held,
nationerna	the nations,nations,
blommor	flowers,
scott	scott,
kvinnors	women's,
aktiviteter	activities,
radion	radio,
vietnamkriget	the vietnam war,vietnam war,
kromosomer	chromosomes,
humör	mood,
alla	all,
protestanter	protestants,
caesars	caesars,
miljön	the environment,
termen	the term,
stadshus	town hall,
samhällets	of society,
tävlingar	competitions,
producerad	produced,
inledande	initial,
produceras	produced,
grekisk	greek,
producerat	produced,
introducerade	introduced,
producerade	produced,
olycka	accident,
budskap	message,
målning	painting,
graviditet	pregnancy,
blodet	the blood,
genom	through,
enstaka	occasional,
england	england,
populärt	popular,
populära	popular,
blues	blues,
förespråkade	advocated,
kretsen	the order,
finner	finds,
uppfördes	was constructed,
kopplad	connected,
garvey	garvey,
norska	norwegian,
uppstått	arisen,
sammanfattning	summary,
besökte	visited,
kopplat	connected,
ingående	enter into,
medel	middle,
sparken	gets fired,
alltmer	increasingly,more and more,
stjärnor	stars,
driver	drive,
både	both,
kostade	cost,
ålands	Åland island's,
poeten	the poet,
teknologi	technology,
turistmål	tourist attraction,
gatorna	the streets,
skolan	school,
nivåer	levels,
besök	visit,
uppenbarelse	apparition,
bidragit	contributed,
relationer	relations,
skiftande	shifting,
spekulationer	speculations,
såg	saw,
gemensamma	common,
liknas	compared to,
sår	wound,
besläktat	related,
läggas	laid,
tappade	lost,
zeus	zeus,
borgmästare	mayor,
moder	mother,
grace	grace,
obama	obama,
återkom	returned,
marknadsekonomi	market economy,
nikolaj	nikolaj,
avslutade	ended,finished,
inkluderar	includes,
generationen	the generation,
inkluderat	including,
generationer	generations,
finansiera	finance,
framåt	forward,forth,
varianten	version,
norstedts	norstedt's,
kongokinshasa	democratic republic of the congo,
varianter	diversities,
vinterspelen	winter games,
sträcker	stretches,
sydostasien	south east asia,
brooklyn	brooklyn,
plan	level,
längtan	longing,
arter	species,
utsattes	subjected,
cover	cover,
kanalen	the channel,channel,
kanaler	channels,
monarki	monarchy,
förklaringen	the explanation,
mesopotamien	mesopotamia,
golf	golf,
pengarna	the money,
presidentens	the presidents,
detalj	detail,
karaktär	character,
falskt	false,
framgångar	successes,success,
existensen	existence,
wayne	wayne,
betydelsen	the meaning,
jämfört	compared,
kontor	office,
gratis	free,
evolutionen	the evolution,
tekniken	techinque,the technology,
tekniker	technician,
föll	fell,
victoriasjön	lake victoria,
tanken	idea,
ledare	leader,
bytet	the exchange,
populärmusik	popular music,
kill	kill,
någon	someone,
kriterier	criteria,
ser	sees,
förhöjd	enhanced,
sex	six,
lyckas	succeed,
järnväg	railway,
något	something,any,
sorters	kinds of,
påverkat	influenced,
guinea	guinea,
fission	fission,
stärkelse	starch,
alqaida	al-qaida,al-qaeda,
rita	draw,
europa	europe,
giftermål	marrige,marriage,
medveten	aware,
avvikelser	deviations,
medvetet	consciously,
stadsdel	district,
utkom	issued,
forskare	scientists,
bästa	best,
medicinering	medication,
förändring	change,
bäste	best,
messias	messiah,
stå	stand,
kopia	copy,
transeuropeiska	transeuropean,
bell	bell,
krisen	the crisis,
allierade	allied,
decennium	decade,
koalition	coalition,
väntade	waited,
tillväxt	growth,
idén	the idea,idea,
föranledde	brought about,
beskrevs	was described,
skönhet	beauty,
östafrika	east africa,
fira	celebrate,
hovrätten	the court of appeal,
fritz	fritz,
uppleva	experience,
systematik	systematic,
framträder	appear,
projekt	project,
budget	budget,
guldbollen	guldbollen,
bestående	comprising,lasting,
brottslighet	criminality,
pressen	the pres,
von	von,
titanic	titanic,
strävar	strives,
lokaler	place,
korruptionsindex	corruption index,
kritiker	critics,
barney	barney,
möjlighet	oppertunity,possibility,
skalet	shell,
barnen	children,
kritiken	the criticism,
laddning	charge,
centrum	center,
snarare	rather,
republiken	the republic of,the republic,
debatten	the debate,
kring	around,
avlägsna	remove,
euro	euro,
normala	normal,
krigsmakt	military power,
person	person,
kontakter	contact,contacts,
nacka	nacka,
tunnelbana	subway,
stränder	beaches,
släppas	be released,
stockholms	stockholm's,
finansiella	financial,
kontakten	the contact,
mandat	mandate,
fascistiska	fascistic,
festivalen	the festival,
nordväst	north west,
festivaler	festivals,
jönssonligan	jönssonligan,
stundom	somtimes,
format	shaped,
teologiska	theological,
melker	melker,
avvisar	reject,
ivar	ivar,
skarp	sharp,
utlösa	trigger,
informationen	the information,
ivan	ivan,
tidigt	early,
lenin	lenin,
saknar	lacks,
saknas	missing,
användbar	useful,
läste	read,
brasilianska	brasilian,
trafiken	the traffic,
turnerade	toured,
religion	religion,
riksförbundet	national association,
säger	says,
nybildade	newly formed,
tåg	trains,
styrelsen	the board,
vagnar	carriges,
plocka	pick,
engelska	english,
bokstav	letter,
engelske	english,
by	village,
ideologin	the ideology,
bosättningar	settlements,
soldaterna	the soldiers,
dagligen	daily,
gemenskaperna	communities,community,
papper	paper,
inte	not,
clinton	clinton,
efterföljande	subsequent,
spridas	spread,
kraven	the demands,
popsångare	pop singer,
uppkallad	named,
seger	victory,
veckor	weeks,
utbröt	erupted,broke out,
knuten	tied to,knot,
fattigdom	poverty,
förbindelse	connection,
européerna	europeans,
poster	positions,
rörlighet	movement,
betyda	mean,
begreppen	the concepts,
begreppet	concept,
atom	atom,
kritisk	critical,
lovade	promised,
lina	lina,
fader	father,
cia	cia,
ut	out,
up	up,
ur	out,
uk	uk,
testamente	will,
öland	öland,
nämner	mentions,
pernilla	pernilla,
utbyggt	built,
personlighetsstörning	personality disorder,
gestalter	figures,
räkna	count,
edwards	edward's,
innehåller	contains,
nordafrika	north africa,
matematiker	mathematician,
besegra	defeat,
dominerades	was dominated,
förstå	understand,
radikala	radical,
djurgårdens	djurgården's,
regissör	director,
riskerar	risks,
springsteen	springsteen,
radikalt	radically,
slås	is hit,
hells	hells,
land	country,
passagerarna	passengers,the passengers,
uppträdande	performance,conduct,
symtom	symptom,
produkt	product,
härstammar	stems,
texten	the text,
inspelning	recording,
persbrandt	persbrandt,
släpptes	was released,
alltför	all too,way too,
bakåt	backwards,
turkisk	turkish,
dyraste	most expensive,
hamnar	lands,
hamnat	ended up,
dickinson	dickinson,
märken	sign,
hustru	wife,
palestinier	palestinians,
kommunistiska	communistic,
drogen	the drug,
tillhörande	belonging to,
påverka	influence,
eva	eva,
jobbet	the job,
romerska	roman,
överlevt	survived,
opinionen	opinion,
agera	act,
leonardo	leonardo,
bolsjevikerna	the bolsheviks,
natur	nature,
förkortningar	abbreviations,
pris	price,
antog	adopted,
expressen	expressen,
indiens	indias,
suveräna	terrific,
möjliggör	enables,
birk	birk,
indian	indian,
ledande	leading,
led	suffered,
lee	lee,
lyckades	succeeded,
leo	leo,
begravd	buried,
motorvägarna	the highways,
casino	casino,
teoretisk	theoretical,
anländer	arrives,
tillkom	resided,
högsta	highest,
opinion	opinion,
huvudvärk	headache,
förlora	lose,
oxenstierna	the oxenstierna,
mening	sentence,
anatolien	anatolia,
varmare	warmer,
rico	rico,
hemlig	secret,
elever	students,
godkänna	approve,
klaviatur	keyboard,
orkester	orchestra,
siffror	numbers,
författning	constitution,
samspel	teamwork,
villor	villas,
lokalt	locally,
lokala	local,
process	process,
etta	number one,first,
high	high,
professor	professor,
syre	oxygen,
sydöstra	south east,
frågor	questions,
saknade	missed,
delad	divided,
västerbottens	västerbottens,
delas	shared,
delar	parts,
sydvästra	southwest,
kriminella	criminal,
amerika	america,
djurens	the animals,
profeten	the prophet,
regeringsmakten	government power,
väckt	awaken,
reagans	reagan's,
or	or,
lundgren	lundgren,
nancy	nancy,
kvinnliga	female,
byggnadsverk	building,
borde	should,
handboll	handball,
hårdast	the hardest,
universiteten	the universities,
frånvaro	absence,
hunnit	had time to,
universitetet	the university,
solvinden	the solar wind,
övergrepp	assault,
eliten	the elite,
uppdelat	split,
tecknet	the sign,
uppdelad	divided,split,
beståndsdelar	elements,
ovanlig	uncommon,
bekant	acquaintance,
hemmaplan	home,
dock	nevertheless,
indikerar	indicates,
rotation	rotation,
sönder	broken,
peking	beijing,
välfärd	wealth,
fortsätta	continue,
smallwood	smallwood,
fördrevs	was banished,
överföras	transferred,
astronomer	astronomers,
intresset	the interest,
banan	banana,
matrix	matrix,
enskilda	individual,
kapitalismens	capitalism,capitalism's,
bekräftades	was confirmed,
undertecknades	signed,
redskap	device,
egenskaperna	the qualities,
påverkats	affected,
förts	brought,
tempererat	temperate,
dubbel	double,
våldsam	violent,
krävs	needs,
david	david,
blanda	mix,
krets	circuit,
helst	rather,
hussein	hussein,
skillnad	difference,
åring	year old,years,
jesus	jesus,
användningsområden	possible use,applications,
nordkoreanska	north korean,
värdefulla	valueable,
festival	festival,
system	system,
tränga	cut in,
teatern	the theater,
blivit	become,
utbyggnad	development,expansion,
haven	the seas,
hampa	hemp,
roberto	roberto,
grundarna	founders,
vecka	week,
jonatan	jonatan,
räcker	enough,
användaren	the user,
filosofin	philosophy,the philosophy,
skick	state,
linda	linda,
viss	certain,
slutsatsen	the conclusion,
nät	web,
minoritet	minority,
slovakien	slovakia,
vardagen	the weekday,
napoleons	napoleon's,
flyga	fly,
medan	while,
framgår	will be seen,
synliga	visible,
våren	the spring,
bokstaven	the letter,
närmade	approached,
brev	letter,
beteende	behaviour,
uppdelade	divided,
manchester	manchester,
hopp	hopes,
östfronten	the east front,
viktor	viktor,
religionens	religion's,
jah	jah,
jag	i,
ilska	anger,
abba	abba,
parlamentet	the parlament,
lägger	put,lies,
fotbollsspelare	football player,
generalen	the general,
bonde	farmer,
britterna	the brits,
h	h,
rowling	rowling,
effekterna	effects,
iranska	iranian,
rymmer	holds,
guvernör	governor,
myndigheterna	the authorities,
debuterade	debuted,
michail	michail,
priser	prizes,
priset	the prize,
lämplig	suitable,
minns	remembers,remember,
vietnams	vietnam's,
författarskap	the writer,authorship,
upprättandet	establishment,
längst	longest,
sjönk	sunk,
balansen	balance,the balance,
bolivias	bolivia's,
enda	only,
bilar	cars,
förklaringar	explanations,
kedjor	chains,
islamiska	islamic,
marknaden	the market,
figuren	the character,
tycker	thinks,
egypten	egypt,
ogillade	disliked,
utövade	exercised,
tätbefolkade	densely populated,
ekvatorn	the equator,
botten	bottom,
dör	dies,
malcolm	malcolm,
mengele	mengele,
sannolikhet	probability,
stabila	stable,
öst	east,
dök	dove,turned,
växa	grow,
keltiska	celtic,
företaget	the company,
moraliskt	morally,
överallt	everywhere,
växt	plant,
genetik	genetics,
louisiana	louisiana,
företagen	the companies,
bilmärke	car make,
molekyler	molecules,
lp	lp,
undervisningen	the education,
atlanta	atlanta,
mandatperiod	term of office,
erhöll	recieved,
rikets	the realms,
demokrati	democracy,
aktivitet	activity,
vd	ceo,
ondskan	the evil,
förlopp	process,developments,
omnämns	is mentioned,
vi	we,
kurdistan	kurdistan,
vm	world championship,
flickor	girls,
skapare	creator,
föreligger	exist,
sitt	its,
referenser	references,
känt	known,
juan	juan,
medeltida	medival,
huden	skin,
romance	romance,
känd	known,famous,
terrorism	terrorism,
flesta	most,
columbia	colombia,
sade	said,
framförde	presented,
homosexuell	homosexual,
anfield	anfield,
ikea	ikea,
diabetes	diabetes,
lupus	lupus,
mänskligt	human,
väger	weighs,weight,
vägen	the road,
mänskliga	human,
uno	uno,
versaillesfreden	treaty of versailles,
paus	paus,
aktuell	current,
renässansen	the renaissance,
paul	paul,
flest	the most,
guds	god's,
förknippas	associated to,
planeter	planets,
frågan	the question,
englands	england's,
planeten	the planet,
filmens	the film's,
förknippad	associated,
motorvägen	highway,
gul	yellow,
dess	its,
arbetarklassen	working class,the working class,
tillverkning	production,
pressas	pressed,
lät	had,
emma	emma,
lär	teach,
vallhund	herding dog,
stadsbild	cityscape,
amazonas	the amazon rainforest,
symptomen	the symptoms,
högskolan	university,
flotta	fleet,
miniatyr|	miniature,
anarkismen	the anarkism,
lägsta	lowest,
transport	transportation,
skriftliga	written,
sällskapet	the company,
toppar	tops,
sålt	sold,
naturlig	natural,
ateist	atheist,
svaga	weak,
biologi	biology,
överlevnad	survival,
östberlin	east berlin,
svagt	weak,
gandalf	gandalf,
smärta	pain,
vargen	the wolf,
användande	use,
kontinenten	the continent,
blodiga	bloody,
angeles	angeles,
upplösningen	disbandment,
planetens	the planets,
kristus	christ,
mera	more,
lycka	happiness,
peters	peters,
skola	school,
överbefälhavare	commander-in-chief,
tina	thaw,
förra	last,
apollo	apollo,
socialistiska	socialistic,
ledamöter	commissioners,
ruset	the fuddle,
stormakt	great power,
monument	monument,
inrättades	established,were implemented,
vanligen	usually,
leukemi	leukemia,
separerade	separated,
särskild	particular,
vitryssland	belarus,
månader	months,
öga	eye,
distinkta	distinct,
särskilt	especially,
modernistiska	modernistic,
övergång	transition,
francisco	fransisco,
uttalade	spoke,
tider	times,
förhandlingar	negotiations,
bröt	broke,
tiden	time,
inspiration	inspiration,
syskon	siblings,
sänker	sinks,
mineraler	minerals,
provinser	provinces,
kommersiell	commercial,
nederländska	dutch,
brevet	the letter,letter,
näsan	the nose,
tätort	conurbation,
preussen	prussia,
bäst	best,
atlanten	the atlantic ocean,
bibel	bilble,
spel	game,
edward	edward,
nervsystemet	the nervous system,
ren	clean,
konsekvens	consequence,
mördade	murdered,
konsekvent	consistent,
golvet	the floor,
främste	premier,
jacob	jacob,
skolor	schools,
innefattar	includes,
slutliga	evenutal,
estland	estland,
jamaica	jamaica,
ständerna	the cities,
galax	galaxy,
horn	horns,
italiens	italy's,
kraftfull	forceful,
tolv	twelve,
bidrag	contribution,
cyklar	bicycles,
bidrar	contributes,
petra	petra,
musikalen	the musical,
räddar	saves,
bortgång	passing,
pluto	pluto,
rapporterar	reports,
begått	committed,
olsson	olsson,
studeras	is studied,
sidan	side,
interstellära	interstellar,
regerande	ruling,
förblir	remains,
stoft	dust,
träda	emerge,fallow,
placerades	placed,
diameter	diameter,
faktiskt	actually,
bro	bridge,
total	total,
bra	good,
stått	stood,
sarah	sarah,
regenter	monarchs,
debutalbumet	the debut-album,
indiana	indiana,
nederlag	defeat,
supportrar	supporters,
riksväg	national highway,
nku	nku,
lissabonfördraget	treaty of lisbon,
friheten	liberty,
fascismen	the fascism,fascism,
era	yours,
specialiserade	specialized,
vietnamesiska	vietnamese,
ekonomiskt	economical,
in	in,
indien	india,
indier	indians,
enhet	unit,entity,
valborg	valborg,
utlandet	abroad,
gotlands	gotland's,
ansluter	connects,
firas	celebrate,
firar	celebrates,
gillar	likes,
sammansatt	composed,
biografer	movie theaters,
neutralt	neutral,
lag	law,
biografen	movie theater,
orden	the words,
medlemsstat	member state,
lämningar	remnants,
livets	life's,
över	over,
office	office,
sovjet	soviet,
exempel	example,
ramadan	ramadan,
söderut	south,
blandning	mixture,
japan	japan,
straff	punishments,
endast	merely,
lagets	the team's,
vanligtvis	usually,
band	band,
fredsbevarande	peacekeeping,
bana	course,
they	they,
spelningen	the gig,
bank	bank,
huvudartikel	main article,
dåliga	bad,
diskuteras	discussed,
knutpunkt	hub,
carlos	carlos,
erbjöd	offered,
germanska	germanian,
inflytandet	the influence,
kejserliga	imperially,
asteroidbältet	the asteroid belt,
trafik	traffic,
bruttonationalprodukt	bnp,
oskar	oskar,
vete	wheat,
klimatet	climate,
nationalistiska	nationalistic,
standard	standard,
tillbaka	back,
berör	affect,concerns,
väldiga	immense,vast,
professionell	professional,
förmågan	the ability,
önskar	wish,
statskupp	coup,
ingmar	ingmar,
kantonerna	cantons,
begränsas	limited,
begränsar	limits,
ingen	no,
begränsat	limited,
förklarade	explained,
förklara	explain,
växthusgaser	greenhouse gas,
inget	no,
john	john,
medborgare	citizens,
antisemitismen	anti-semitism,
äter	eat,eats,
militärt	military,
albert	albert,
kvarvarande	remaining,
persson	persson,
trupp	troops,troop,
finska	finnish,
roms	romes,
symboliserar	symbolizes,
sonen	the son,
används	use,
byggts	built,
minut	minute,
årens	the year's,
skolorna	the schools,
mannen	the man,
onani	masturbation,
omvandling	transformation,
kallades	was called,summoned,
småningom	eventually,
kalendern	calender,
magnus	magnus,
sjukvård	healthcare,
aftonbladet	aftonbladet,
lades	put,
anatomi	anatomy,
närvaro	attendance,
historisk	historical,
verkar	seems,
flygplatser	airports,
bruce	bruce,
utställning	exhibition,
fjädrar	feathers,
flygplatsen	the airport,
aminosyra	amino acid,
ägda	owned,
ägde	owned,
bortom	beyond,
läran	the teaching,
evigt	forever,
misslyckade	failed,
förväxla	mistake,
effekten	the effect,
mitten	middle,
hinduiska	hindu,
madeira	madeira,
tilläts	was allowed,
senare	later,
fortplantning	reproduction,
rankning	ranking,
sättet	manner,
 kilometer	kilometer,
sätter	place,puts,
kejsar	emperor,
inställning	attitude,
målvakt	goalee,
kontinuerlig	continuous,
dj	dj,
de	the,
sverigedemokraterna	sweden democrats,
stalins	stalins,
orolig	worried,
du	you,
dr	doctor,
offret	the victim,
runt	around,
spridningen	the spread,
konst	art,
tyngre	heavier,
fågelarter	species of bird,
lasse	lasse,
libanon	lebanon,
kurdiska	kurdish,
vanlig	ordinary,
utförd	completed,performed,
treenigheten	the trinity,
historiens	historys,
sexuell	sexual,
djuret	the animal,
fångenskap	captivity,
materialet	the material,material,
smaken	the flavour,
we	we,
intog	seized,occupied,
miljö	environment,
jämförelse	comparison,
huvudsakligen	primarily,
garanterar	ensures,guarantees,
kännetecknas	is characterized,
brad	brad,
målningen	the painting,
graviditeten	the pregnancy,
kännetecken	distinction,
thierry	thierry,
fångar	prisoners,
chrusjtjov	chrusjtjov,
genomför	implement,
tony	tony,
smith	smith,
japans	japans,
patienten	the patient,
framträdande	apperance,
huvud	head,
hitlers	hitlers,
patienter	patients,
attacken	the attack,
attacker	assaults,
fest	party,
juridik	law,
drottningen	the queen,
frekvens	frequency,
vagn	carrige,
johansson	johansson,
påstådda	alleged,
kupp	kupp,
nordöstra	nordeastern,
spanjorerna	the spaniards,
have	have,
moldavien	moldova,
deltagarna	participants,
påverkades	was affected by,
själva	self,
våg	road,
patent	patent,
utgivna	published,
ersattes	was replaced by,
andelen	the share,the proportion,
raid	raid,
hann	reached,
balkan	the balkans,
sexualitet	sexuality,
delstaten	the state,
hans	his,
bilen	the car,
koncentrerad	concentrated,
aspekter	aspects,
rörelsen	movement,
somliga	some,
styrkorna	forces,
mamma	mother,
röd	red,
gärningsmannen	culprit,
newton	newton,
kall	cold,
nästan	almost,
kroppens	the body's,the bodies,
kalender	calender,
swahili	swahilli,
så	so,
distributioner	distributions,
havets	the seas,
kritiska	critical,
plasma	plasma,
född	born,
maya	maya,
återgick	returned,returning,
skadorna	damages,
arab	arab,
fusion	fusion,
indianer	indians,
uppträdde	perform,
everton	everton,
engelskans	english,
hepatit	heptatitis,
årlig	yearly,
indelning	the subdivision,
indelningen	division,
samfund	order,
gandhi	gandhi,
transkription	transcript,
sixx	sixx,
bort	away,
presidentvalet	presidential election,
borg	tower,castle,
bord	table,
humor	humour,
serbiens	serbias,
siffran	number,
stadsdelarna	districts,
vägar	roads,
bevara	preserve,
vunnit	won,
juryns	the jury's,
jacques	jacques,
återfinns	is rediscovered,
karlsson	karlsson,
kommittén	the committee,
efternamn	lastname,
gemenskapen	the collective,community,
way	väg,
war	war,
etablerat	established,
skiljas	separate,
motorvägar	highways,
inträffar	occur,
partiledare	party leader,
emil	emil,
reser	travels,
studierna	the studies,
litterär	literary,
långvarig	long,
träning	training,
erövra	conquer,
engagerade	engaged,
utomlands	abroad,
xiis	xii,
efter	after,
bilderna	the pictures,
empati	empathy,
toppen	the top,
arkitekten	the architect,
förmåga	ability,
janukovytj	janukovytj,
knäppupp	knäppup,knäppupp,
arkitekter	architects,
test	test,
götaland	götaland,
konservatism	conservatism,
mött	met,
femton	fifteen,
reglerar	regulates,
regleras	is regulated,
omgivande	surrounding,surounding,
rätten	the court,
bergmans	bergman's,bergmans,
uppfanns	was invented,invented,
global	global,
datum	date,
redaktör	editor,
lider	suffers,
utkämpades	fought,
afrikaner	africans,
rådet	council,
råder	advises,
ätten	the dynasty,
vänder	turn,
division	division,
uttrycka	express,
lättare	easier,
hannar	males,
uttryckt	expressed,
enskilt	individually,
konstnärlig	artistic,
datorspel	video game,
levnadsstandard	standard of living,
frigörs	is released,
litterära	literal,
revolution	revolution,
alfa	alpha,
engagerad	engaged,
invandrade	immigrated,immigrant,
sköttes	operated,
motsatte	opposed,
stimulera	stimulate,
motsatta	opposite,
ungdomar	youths,
ingick	were included,
kosmiska	the cosmic,
fastigheter	real estates,
utspelar	takes place,set,
gener	genes,
marxismen	marxism,
kärlek	love,
påstår	claims,asserts,
genen	the gene,
oerhört	tremendously,
antarktiska	antarctic,
sistnämnda	later,
kemi	chemistry,
franklin	franklin,
ponny	pony,
vinnare	winner,
ekr	ekr,
dåtidens	past times,that time,
vapnet	the weapon,
spridit	spread,
vapnen	the weapons,
förteckning	listing,
kärnkraftverk	nuclear power plant,
presenterar	presents,present,
upprättade	established,
stabilitet	stability,
regel	rule,
omvärlden	surrounding world,
fransmännen	the french,
snabbt	quickly,
målvakten	the goalkeeper,
ämnena	the elements,
närmar	close in,closing,
varför	why,
norrköpings	norrköpings,
snabba	rapid,
löner	salaries,
ibm	ibm,
ibn	ibn,
interaktion	the interaction,interaction,
frukt	fruit,
erbjuder	offers,
några	a few,
december	december,
nobels	nobel's,
gentemot	towards,against,
abort	abortion,
genomgått	experienced,
ligan	league,
pojke	boy,
betydelse	significance,
kopplingar	connections,
perserna	the persians,
göteborgs	gothenburgs,
ungern	hungaria,
stöds	is supported,
flyttas	moved,
flyttar	move,
kurs	course,
rekordet	the record,
maktens	the powers,the power's,
landshövding	county governor,
ganska	quite,
ättlingar	descendants,
magnetfält	magnetic field,
generalguvernören	general governor,
fält	field,
skabb	scabies,
levde	lived,
utnämndes	was declared,
därifrån	from there,
bergskedjan	the mountain group,
nominerades	was nominated,nominated,
hals	throat,
halt	stop,
varar	lasts,
nog	enough,
författarna	writers,
förvaras	is stored,
komponenter	components,
terrorismen	the terrorism,
now	now,
frihet	freedom,
språk	language,
antyder	indicates,
stockholm	stockholm,
januari	january,
drog	draw,
em	european championship,
sektorn	the sector,
citat	quote,
ed	ed,
utbrett	wide,
strålningen	radiation,
eu	eu,
et	et,
kant	kant,
fuglesang	fuglesang,
ep	ep,
er	you,
album	album,
teorier	theories,
återkommande	recurring,
stallone	stallone,
koffein	caffein,
carl	carl,
sven	sven,
domen	judgment,
allmänheten	general public,
xi	xi,
derivatan	the derivative,
bergqvist	bergqvist,
omtvistat	disputed,
desmond	desmond,
sheen	sheen,
satsningar	investments,
färre	less,
fascisterna	fascists,
television	television,
europeisk	european,
sidorna	the pages,pages,
ändrades	changed,
kloster	monastery,
grundad	founded,
craig	craig,
statsminister	prime minister,
kairo	cairo,
grundar	bases,
anges	is put at,
hjälp	help,
hör	hears,
fortsatta	continued,
etiopiska	ethiopian,etiopian,
bönor	beans,
hög	high,
skäl	reasons,
numera	now,
bön	prayer,
bekostnad	expense,
dvärgar	dwarfs,
glödlampor	light bulbs,
america	america,
på	on,
michelle	michelle,
lyfter	lifts,
norrmän	norwegians,
nordligaste	northern,
runda	round,
orsaka	cause,
abraham	abraham,
skapats	was created,
kyrkorna	the churches,
marocko	marocco,
teori	theory,
perfekt	perfect,
rötter	roots,
huskvarna	huskvarna,
sierra	sierra,
definierade	defined,
uppståndelse	resurrection,
helgdagar	holidays,
riddare	knight,
samuel	samuel,
mission	mission,
ambitioner	ambitions,
folkomröstning	referendum,
facupen	fa-cup,
bushadministrationen	the bush administration,
storstäder	metropolises,
sport	athletics,sport,
katastrofer	catastrophes,
depressionen	the depression,
konstaterade	established,
ladin	ladin,
depressioner	recessions,
israels	israel's,
import	import,
kommunismens	the communisms,
katastrofen	the catastrophy,
yta	surface,
personlighet	personality,
utgivningen	the publication,
rike	kingdom,
utgavs	was published,
samtal	call,
warhol	warhol,
rika	rich,
kristinas	kristina's,
feminismen	feminism,
ståndpunkt	standpoint,
nils	nils,
placerar	places,
placeras	placed,
avskaffande	abolition,
dömande	judging,
bomull	cotton,
östtyska	east german,
handlande	action,
långfilm	feature film,
oliver	olives,
lyssnade	listened,
oden	oden,
knappt	barely,
dräkt	costume,
observera	observe,
utförda	made,performed,
elvis	elvis,
funnits	been,
ytan	area,
uefacupen	the uefa champions league,
prinsessan	the princess,
polens	polands,
ordningen	the order,order,
ansikte	face,
tjeckien	czech republic,the czech republic,
eran	era,
beläget	base,
inslag	elements,
finanskrisen	the financial crisis,
behandlade	treated,
kvarter	quarter,block,
kenya	kenya,
helium	helium,
infödda	natives,
slaget	the strike,
programvara	software,
långa	long,
homosexualitet	homosexuality,
pesten	the plague,
lite	little,
speciella	special,
offensiven	offensive,
skivbolaget	record label,
acdc	ac/dc,
omfattande	large,
målningar	paintings,
omfattas	comprise,
omgående	immediate,
tradition	tradition,
fredspris	peace prize,
erkänd	acknowledged,
flaggor	flags,
mynning	outfall,mouth,
forskarna	the scientists,
skandinaviska	scandinavic,
framgången	the success,
eleverna	the pupils,the students,
lagerkvist	lagerkvist,
nazismen	nazism,
euron	the euro,
ca	cirka,
lade	laid,
slöts	signed,
irland	ireland,
passiv	passive,
stund	while,
östergötland	Östergötland,
selma	selma,
amy	amy,
symbolisk	symbolic,
strävan	the quest,
skilda	separate,
varandra	each other,
eddie	eddie,
lågt	low,
präglades	imprinted,
slår	beats,
användbara	usable,
sålts	sold,
kategoripersoner	category of persons,
berodde	depended,
innebörden	the significance,
utskott	organ,
bestämt	decided,
nsdap	nsdap,
jussi	jussi,
bestäms	is decided,
kaffet	the coffee,
francis	francis,
ideologi	ideology,
palme	palme,
central	central,
sri	sri,
bidragen	contributions,
efterkrigstiden	the post-war period,
kapten	captain,
klassiker	classic,
karriär	career,
area	area,
specifikt	specifically,
stark	strong,
start	start,
anställd	hired,
specifika	specific,
likväl	nevertheless,still,
gånger	times,
fastställa	determine,confirm,
hawking	hawking,
guillou	guillou,
wailers	wailers,
sämsta	worst,
gången	time,
traditionerna	the traditions,
expeditionen	the expidition,
minne	memory,
freddy	freddy,
miguel	miguel,
expeditioner	expeditions,
kostar	costs,
godkände	approved,
knut	knut,knot,
evenemang	event,
nere	down,
mongoliet	mongolia,
upphovsman	author,creator,
tänderna	teeh,
drift	drift,
massachusetts	massachusetts,
röda	red,
skuggan	the shadow,
tjänare	servant,
morgonen	the morning,
olympiastadion	olympa stadium,
eriksson	eriksson,
beskrivningar	descriptions,
energikälla	energy source,
öknen	the desert,desert,
antoinette	antoinette,
griffin	griffin,
påbörjades	was started,
lämpligt	suitable,
skiljer	differs,
får	can,
verk	work,
tredje	third,
heaven	heaven,
sverige	sweden,
behöver	need,
louis	louis,
resan	the trip,
koranen	the quran,
rasism	racism,
magdalena	magdalena,
fåglarnas	the birds',
egendom	property,
orgasm	orgasm,
markerade	marked,
trupper	troops,
utåt	outwardly,
höja	raise,
tvskådespelare	tv actor,
bedrev	managed,
bernhard	bernhard,
misstänkta	suspected,
förbjudet	prohibited,
irak	iraq,
genomförde	carried out,
kronor	kronor,
observeras	observed,
uttalat	outspoken,
lämna	leave,
uttalas	pronounced,
arena	arena,
vår	spring,
krigen	wars,
externa	external,
minst	at least,
boxning	boxing,
sagor	fairytales,
kriget	the war,
hoppades	hoped,
perspektiv	perspective,
då	then,
nazityskland	nazi germany,
grunda	found,
kritiserat	criticised,
nukleotider	nucleotides,nucleotide,
familj	family,
avsedd	intended,
avgör	decides,
arrangemang	arrangement,
taket	the roof,
bolagets	the corporation's,
representeras	represented,
expansionen	the expansion,
ryssland	russia,
reptiler	reptiles,
utökat	extended,
blodtryck	blood pressure,
latinamerikanska	latin american,
räknat	counted,
räknar	counts,
lagstiftande	legislating,
ständigt	always,
gazaremsan	the gaza strip,
ombord	onboard,
livslängd	life expectancy,
feministiska	feminist,
gälla	be valid,
serber	serbs,
linköping	linköping,
reidars	reidars,
utför	perform,
betraktades	regarded,
fastän	although,
fd	ex,
samarbeten	collaborations,
fn	the un,
vattenkraft	hydroelectric power,
kostnaden	cost,
byggandet	the building,
enzymer	enzymes,
segrar	victories,
skiljs	separate,
kostnader	expenses,
dream	dream,
nämnts	mentioned,
tillgångar	assets,
helt	totally,
tornet	the tower,
tornen	towers,
hela	entire,
hell	hell,
kombinerade	combined,
hundratusentals	hundreds of thousands,
paulo	paulo,
hendrix	hendrix,
systems	systems,
österrikes	austria's,austrias,
musikalisk	musical,
bytte	swapped,
elden	the fire,
konstitutionella	constitutional,
greps	was arrested,
dyrt	dearly,
petter	petter,
fullt	completely,
fulla	complete,
skrivit	written,
kontinentens	the continents,
ifk	ifk,
etnisk	ethnic,
positionen	the position,
rättvisa	justice,
försäljning	sales,sale,
aktörer	players,
robert	robert,
bodde	lived,
lungorna	the lungs,
stödet	the support,
stöder	supporting,
utredningen	the investigation,
heroin	heroine,
vasas	vasas,vasa's,
svarade	answered,
skilja	seperate,
underhåll	allowance,
ytterligare	additional,
sänder	broadcast,transmits,
sändes	was sent,
etiska	ehtical,
arsenal	arsenal,
minoritetsspråk	minority language,
synes	seems to,appears,
miss	miss,
rygg	back,
deltagare	contestant,
kongresspartiet	indian national congress,
station	station,
parlamentsvalet	parliament election,
nigeria	nigeria,
kallar	calls,
brittiska	british,
luminositet	luminosity,
läsa	read,
åkte	relegated,
representera	represent,
förnuftet	reason,
brittiskt	british,
tvungen	forced,
växterna	plants,
stora	big,
långsamt	slowly,
einsteins	einsteins,
andersson	andersson,
värden	values,
värdet	the value,
gren	branch,
charlotte	charlotte,
bestämdes	was determined,
teslas	tesla's,
genomgripande	good,
tvärtom	on the contrary,contrary to,
nominerad	nominated,
militär	military,
demokratin	the democracy,
liberalismen	the liberalism,
lik	similar,alike,
liv	life,
herre	lord,
avseenden	regard,
måne	moon,
mexiko	mexico,
världsarvslista	world heritage list,
freddie	freddie,
kap	chapter,
utgör	constitutes,
himlakroppar	celestial bodies,
södra	south,
polacker	poles,
räknade	counted,
recensioner	reviews,
två	two,
ingenting	nothing,
deltar	participates,
möjligen	possibly,
counterstrike	counterstrike,
muslimsk	muslim,
justice	justice,
humanistiska	humanistic,
åländska	Åland swedish,
ikon	icon,
ingå	be a part,be included in,
avsaknaden	absence,
vilken	which,
ingredienser	ingredients,
västkusten	the west coast,
maurice	maurice,
bakgrund	background,
tidigare	earlier,
ändamål	purpose,
mörkare	darker,
direktör	director,
upphovsrätten	copyright,
pjäser	plays,
löst	solved,
allvar	earnest,
likhet	similar,resemblance,
utsträckning	extent,
revolutionen	the revolution,
länk	link,
lejonet	the lion,
anor	ancestry,
viljan	will,
slavar	slaves,
kyrkliga	religious,from the church,
läsaren	the reader,
uppfylla	satisfy,
betydde	meant,
derivata	derivative,
scientologikyrkan	the church of scientology,church of scientology,
sokrates	socrates,
merparten	most,
minskade	was reduced,
oändligt	infinitely,
gestalt	figure,
walter	walter,
handlingen	the story,
budgeten	the budget,
anthony	anthony,
livet	the life,
delades	split,
socialism	socialism,
hegel	hegel,
läses	is read,
läser	read,are reading,
guide	guide,
slutar	end,
slutat	ended,
uttryckte	expressed,
lagar	laws,
tillfällen	oppertunities,
kombineras	combined,
staffan	staffan,
kombinerat	combined,
ändra	change,
deltagande	participation,
nöd	distress,
kombinerad	combined,
inledde	started,
folkslag	kind of people,
kungahuset	royal house,
anklagats	accused,
kommunicera	communicate,
förlag	magazine,
seglade	sailed,
svealand	svealand,
fatta	make,
kurdisk	kurdish,
flygplan	airplane,
nutid	present,
präglad	marked,characterized,
innersta	innermost,
njurarna	the kidneys,
tortyr	torture,
skal	shell,
fredliga	peaceful,
kallblod	cold blooded,
gänget	the gang,
nikki	nikki,
varuhus	department store,
djup	deep,
huvudort	principal town,
bestå	consists,exist,
producerats	produced,
gör	does,makes,
enklare	simpler,
gitarristen	the guitarist,
immigranter	immigrants,
uppvärmningen	the warm-up,
dylikt	such,
gandhis	gandhi's,
unge	kid,
donna	donna,
begärde	demanded,
mycket	much,
byggnader	buildings,
biträdande	assisting,
pierre	pierre,
våldet	the violence,
economic	economic,
tämligen	fairly,
syndrom	syndrom,
sammanhängande	connective,
skapat	created,
vilda	wild,
skapar	creates,
faktorn	factor,
journalist	journalist,
run	run,
steg	rose,
sten	stone,
mellankrigstiden	interwar years,
naturvetenskapliga	scientific,
socialister	socialists,
benfica	benfica,
bistånd	aid,
führer	fuhrer,
övergick	transended,
efterträdare	successor,
linjer	lines,
edvard	edvard,
länderna	the countries,
ändringar	changes,
ida	ida,
öl	beer,
reaktorer	reactors,
institut	institution,
emellan	between,
föreningen	association,
fokuserade	focused,
visar	shows,
består	exists,
visat	shown,
heritage	heritage,
jonsson	jonsson,
ledamot	representative,
strukturen	the structure,
larry	larry,
strukturer	structures,
drabbats	afflicted,
ute	out,
nyval	re-election,
malin	malin,
trafikerade	frequent,
  km²	square kilometre,
politik	politics,
chelsea	chelsea,
ligacupen	league cup,
bränslen	fuel,
avsåg	meant,
uppfyller	fulfills,
hårdrock	hard rock,
igenom	through,
krigets	the war's,
sjunde	seventh,
berättat	told,
klubbarna	the clubs,
berättar	tells,
berättas	is told,
korn	korn,barley,
rester	remains,
dras	draw,
drar	earn,
drag	move,
mästare	master,
matematiska	mathematical,
resten	the rest,
vindar	winds,
kors	cross,
närmaste	closest,
e	e,
enade	united,
medför	entails,
officerare	officer,
tunga	tongue,
tillfälliga	temporary,
svt	svt,
dvs	i.e.,
bonniers	bonnier's,
höst	autumn,
indiska	indian,
företeelse	phenomenon,
ge	give,
tänker	thinking,
go	go,
träd	tree,
danmark	denmark,
världsrekord	world record,
tillhör	belongs,
flitigt	actively,
ännu	yet,
kommunismen	communism,
ryan	ryan,
utbredning	distrubution,
stift	diocese,
carter	carter,
mussolinis	mussolini's,
honan	the female,
geologiska	geological,
visserligen	certainly,
direkta	direct,
börjar	starts,
träffades	was met,
mussolini	mossolini,
kinas	chinas,
erövringar	conquests,
hansson	hansson,
polen	poland,
gradvis	gradually,
genombrott	breakthrough,
cell	cell,
experiment	experiment,
avancerade	advanced,
gamla	ancient,
utrikespolitiken	the foreign policy,
gamle	old,
offentlig	public,
händelsen	the occurence,
gåva	gift,
eminem	eminem,
ryska	russian,
innebandy	floorball,
västerut	westwards,
ateism	atheism,
kraftig	strong,
uppfinningar	inventions,
avsedda	intended,
italienska	italian,
genetiska	genetic,
personen	the person,
kunde	could,
personer	people,
oktober	october,
mexikanska	mexican,
nordkorea	north korea,
invigningen	the opening,
huxley	huxley,
turkiets	turkey's,
debutalbum	debut album,
befolkningstäthet	population density,
kenny	kenny,
liknade	looked like,
halloween	halloween,
talat	spoke,
talas	is spoken,
talar	speaks,
tåget	the train,
georg	georg,
tågen	the trains,
sovjetunionen	the soviet union,
fälttåg	campaign,
folkmängd	population size,population,
kronprinsen	crown prince,the crown prince,
oroligheter	unrest,
fara	danger,
uttalet	the pronounciation,
svenskar	swedish,
dödlig	mortal,
fart	speed,
utfördes	preformed,
ringde	called,
säljer	sells,
reagerar	reacts,
rörde	had something to do with,touched,was about,
kungliga	royal,
kapital	capital,
högtider	holiday,
fungerade	working,
presidenter	presidents,
förstördes	was destroyed,
någonting	anything,
presidenten	the president,
offentligt	publicly,
verklighet	reality,
belopp	sum,
monarken	the monarch,
insekter	insects,
allting	everything,
naturgas	natural gas,
zagreb	capital of croatia,
ägna	spend,devote,
läror	teachings,
konserter	concerts,
dikt	poem,
intäkterna	the revenues,
miniatyr|px|den	miniature,
hunden	the dog,
kläder	clothes,
räckte	enough,
mode	fashion,
förmågor	capacities,abilities,
modo	modo,
dömdes	was convicted,
föreslogs	was suggested,
illuminati	illuminati,
globe	globe,
skolgång	school attendance,
 procent	percent,
stiger	rises,
osmanerna	ottoman turks,
illa	bad,
flyr	flees,
entertainment	entertainment,
islamisk	islamic,
samarbetar	cooperates,
samarbetat	collaborated,
max	max,
solsystem	solar system,
sedermera	since,
kropp	body,
bilder	pictures,
lida	suffer,
bilden	the image,
förstod	understood,
förbund	union,
kommunala	local,municipal,
banor	paths,line,
densamma	the same,
benämnas	named,
strida	fight,
tillgången	access,
tigrar	tigers,
austin	austin,
riksdagsvalet	parliamentary election,
ursprungsbefolkningen	the native population,
önskemål	requests,
undervisade	taught,
boken	the book,
upphört	ceased,
kulturarv	cultural heritage,
nilsson	nilsson,
hasch	hashish,
styrelseskick	form of government,government,
lista	list,
representerade	represented,
definieras	is defined,defines,
arbetade	worked,
inbördes	intermutual,
israelisk	israeli,
ber	asks,
julian	julian,
bordet	the table,
benämning	term,name,
visor	songs,
förlorades	was lost,
släkt	family,
runorna	the runes,
förblev	remained,
jorge	jorge,
regn	rain,
genomslag	breakthrough,
tyskar	germans,
sändas	be transmitted,
skogar	forests,
långtgående	far-reaching,
platon	platon,
minska	reduce,
församling	congregation,
parken	the park,
hade	had,
basen	became,
radioaktivt	radioactive,
gemensam	common,
härskare	ruler,
varit	been,
överlever	survives,
aspekt	aspect,
psykologin	the psyhology,
boris	boris,
klassiska	classic,
inbördeskrig	civil war,
omloppsbana	orbit,
michigan	michigan,
förbjöd	forbid,
området	the area,
inflytelserika	influential,
klassiskt	classical,
häst	horse,
karriären	the career,
älskade	loved,
gray	gray,
processer	processes,
tillgång	access,
mohammed	mohammed,
grav	grave,
gran	spruce,
influensa	influenza,
också	also,
processen	the process,
vänt	turned,
fru	wife,
sydafrika	south africa,
västindien	west india,
korea	korea,
volvo	volvo,
individens	the individual's,
gotiska	gothic,
staty	statue,
state	state,
företagets	the company's,
ken	ken,
högra	right,
sovjetiska	soviet,sovjet,
benämningen	the name,
jobba	work,
befälet	the command,
nedre	lower,
innanför	inside,
odens	odin's,
vulkaner	volcanos,volcanoes,
nyare	newer,
trädde	come into effect,
varierade	varied,
älskar	loves,
stratton	stratton,
framgångsrikt	successful,
partiklar	particles,
jersey	jersey,
uppsättning	equipment,
fördelar	share,
fördelas	distribute,
torn	tower,
leipzig	liepzig,
genre	genre,
kings	king's,
sammanhang	context,
christer	christer,
liberala	liberal,
äldre	older,
poet	poet,
påminde	reminded,
ämbetsmän	bailies,
kingston	kingston,
vinci	vinci,
spanska	spanish,
spanien	spain,
bär	carryng,berries,here,
strömningar	sentiments,
kanarieöarna	the canary islands,
erbjuda	offer,
könsorganen	the genitals,the reproductive organs,
utgjorde	made up,
avrättades	was executed,
reaktion	reaction,
nordens	the scandinavian countries',
rysslands	russia's,
enkel	simple,
feber	fever,
demo	demo,
rättigheter	rights,
måleri	painting,
alfabetisk	alphabetical,
parti	party,
friidrott	track and field,
campus	campus,
varmed	whereby,
förebyggande	preventive,
växjö	växjö,
flygbolag	airline,
anka	anka,duck,
representerar	represents,
införa	introduce,
nämligen	namely,
infört	introduced,
alperna	the alps,
lagring	storage,
flickan	the girl,
strömmen	the stream,
grenar	branches,
i	in,
theodor	theodor,
onda	evil,
brandenburg	brandenburg,
störta	rush,
sänds	sends,
sofia	sofia,
sofie	sofie,
sände	sent,
vida	wide,
jeff	jeff,
lutning	closing,incline,
nato	nato,
katolska	catholic,
utan	without,
sanning	truth,
vanligare	more common,
historia	history,
historik	history,
klassificering	classification,
loss	unstuck,
norges	norway's,
fernando	fernando,
martin	martin,
page	page,
regeringar	governments,
lager	layer,
kolonierna	colonies,
vardagliga	everyday,
pojkarna	the boys,
homo	homo,
skorpan	crust,
peter	peter,
 km²	kilometres,
jugoslaviska	yugoslavian,
hyser	accomodates,holds,
folkets	the people's,
alliansen	the alliance,
skriften	writings,
broar	bridges,
motsättningar	oppositions,
samlades	collected,
journal	journal,
reza	reza,
expansion	expansion,
halvön	the peninsula,
keramik	ceramics,
freedom	frihet,
beslutade	decided,
göteborg	gothenburg,
troligen	likely,
hävdade	claimed,
mytologi	mythology,
glenn	glenn,
washington	washington,
längsta	longest,
hammarby	hammarby,
museum	museum,
distinkt	distinctive,
neutral	neutral,
ho	ho,
överens	in agreement,
fysik	physics,
pippin	pippin,
förslaget	the suggestion,
bitar	pieces,
farlig	dangerous,
ordbok	dictionary,
ibland	sometimes,
erik	erik,
eric	eric,
diego	diego,
moderaterna	the moderates,
jordbävning	earthquake,
serveras	is served,
vulkaniska	vulcanic,volcanic,
enastående	exceptional,
revolutionära	revolutionary,
stad	city,
resulterade	resulted,
stan	town,
ockupationen	occupation,
hjärnan	the brain,
stam	tribe,
förekomma	occur,
inser	recognize,realizes,
alkohol	alcohol,
blogg	blog,
konsumtion	consumption,
hinner	have time to,
felaktig	incorrect,
andre	other,
buddy	buddy,
likaså	also,
swan	swan,
kommersiellt	commercial,
kulturell	cultural,
kommersiella	commercial,
köpmän	traders,merchants,
gjordes	made,was made,
vasa	vasa,
åstadkomma	create,
upplysningen	the enlightenment,
kända	known,
kände	felt,
examen	exam,
disneys	disneys,
försöka	try,
chokladen	the chocolate,
avståndet	the distance,
okänt	unknown,
sexton	sixteen,
upp	up,
rollfigurer	roll model,
force	force,
förstaplatsen	first place,
dennes	his,
avfall	waste,
neo	neo,
omedelbart	immediately,
kommissionen	the commission,
ned	down,
trodde	thought,
porträtt	portrait,
med	with,
genomföra	perform,
men	but,
drev	drove,
vinden	the wind,
mer	more,
luther	luther,
geografiskt	geographically,
därpå	thereon,
åka	go,
ajax	ajax,
sju	seven,
pilatus	pilatus,
geografiska	geographical,
magnusson	magnusson,
reste	travelled,
efterföljare	following,
rosenberg	rosenberg,
reagan	reagan,
inleddes	began,initiated,
fördelning	distribution,
soldat	soldier,
berättelserna	the stories,
gävle	gävle,
army	army,
provisoriska	provisional,
rockband	rock band,
oscar	oscar,
grundande	founding,
upplevde	experienced,
wikipedias	wikipedias,
köln	köln,
flora	flora,
kapitalistiska	capitalistic,
sundsvall	sundsvall,
kanadas	canada's,
tidskriften	the magazine,
abstrakta	abstract,
världskrigets	the world war's,
förväntade	expected,
talets	the speechs,
konstitutionen	constitution,
tusen	thousands,
tidskrifter	periodicals,
vänster	left,
satt	sat,
nobelstiftelsen	nobel foundation,
bonaparte	bonaparte,
avrättningen	the execution,
trött	tired,
begrepp	concept,
polis	police,
stilla	still,
orsakar	causes,
orsakat	caused,
utomeuropeiska	non-european,
startade	started,
könsorgan	sex organ,
klarar	do,
president	president,
indelat	divided,split,
medföra	result,
indelad	divided,
medfört	led to,
indisk	indian,
borgerliga	conservative,
färdig	done,
förfäder	ancestors,
föreställningen	the concept,
ibrahimović	ibrahimovic,
munnen	the mouth,mouth,
murray	murray,
föreställningar	performances,
helena	helena,
buddhister	budhists,buddhists,
nationell	national,
personal	personal,staff,
förödande	devastating,
irans	iran's,
federationen	federation,
friska	fresh,
förlängning	extension,
infektioner	infections,
startar	begins,
miljon	million,
myntades	coined,was coined,
exakta	exact,
huvudrollen	leading part,
sida	side,
side	side,
kammaren	the chamber,
liga	league,
päls	fur,
enorm	enormous,
medier	media,
håret	the hair,
uppsala	uppsala,
hänvisa	refer,
ihop	together,
talen	years,
gärna	readily,
sluta	end,
återfanns	was rediscovered,
foto	photo,
neutroner	neutrons,
larssons	larsson's,
normer	standards,
nomineringar	nominations,
uppförande	behavior,
folkvalda	elected,
faktum	fact,
iso	iso,
representant	representative,
berömt	praised,
starta	launch,
gå	go,
leddes	was led,
massiv	massive,
objektet	object,
föreslagit	suggested,
vikingatiden	the viking age,
förbi	past,
objekten	the objects,
hollywood	hollywood,
någonstans	somewhere,
åskådare	spectators,
medeltiden	middle ages,
besegrades	defeated,
hundar	dogs,
formell	formal,
kontrast	contrast,
antarktis	antarctica,
street	street,
regissören	director,
troligtvis	probably,
stadsdelen	the district,
låta	let,
mina	mine,
självständigt	independent,
lämnar	leaves,
lämnas	left,
lämnat	left,
skildringar	descriptions,
monetära	monetary,
ulrich	ulrich,
blue	blue,
dessa	these,
bildar	form,
bildas	formed,
norra	northern,
bildat	formed,
luthers	luthers,
diskuterats	discussed,
don	don,
dom	conviction,
dog	died,
slipknot	slipknot,
följande	following,
kristen	christian,
långvariga	long-standing,
införde	introduced,
hjälper	helps,
befälhavare	commander,
droger	drugs,
skyldig	responsible,guilty,
långvarigt	prolonged,long-standing,
odling	cultivation,
krönika	chronicle,
förutsätter	assume,assumes,
monica	monica,
stycke	piece,
meningar	sentences,
dramaten	dramaten,
stop	stop,
stol	chair,
präster	priests,
stod	stood,
bar	bar,
bas	base,
existerat	existed,
förändra	change,
gärningar	deeds,
zonen	the zone,
gunnar	gunnar,
dittills	thus far,
öppnade	opened,
inledningsvis	by way of introduction,
underart	subspecies,
göta	göta,
rörelsens	movements,
smguld	gold medal in the swedish championships,
artikel	article,
armeniska	armenian,
kämpa	fight,
regelbundet	regularly,
isotoper	isotopes,
fns	un's,
regering	the government,
näringslivet	industrial life,
fördraget	the treaty,
fördragen	the compacts,
ung	young,
regelbunden	regular,
obamas	obama's,
rysk	russian,
mellanrum	gap,space,
nationalförsamlingen	national assembly,
hittar	finds,
interna	internal,
omstritt	controversial,
erövrade	conquered,
cyrus	cyrus,
ting	matters,
frisk	healthy,
tillämpa	administer,
betydelsefull	meningful,
igång	start,start up,
utseende	appearance,
sällskapshundar	pet dogs,companion dog,
namnen	names,
mindre	smaller,
förgäves	in vain,
albaner	albanians,
ip	ip,
sushi	sushi,
marco	marco,
sommar	summer,
colosseum	colosseum,
konkurrensen	the competition,
vänstern	western,
make	husband,
bella	bella,
västberlin	west berlin,
kommunistpartiets	the communist partys,the communist party,
roland	roland,
därmed	therefore,
industriell	industrial,
makt	power,
benämningar	terms,
anglosaxiska	anglo-saxon,
atmosfären	the atmosphere,
skickades	was sent,
kim	kim,
nicklas	nicklas,
folkrikaste	most populus,
nedan	below,
vetenskaplig	scientific,
dåvarande	formerly,
värmland	wermlandia,
roma	roma,
grannländer	neighboring countries,
just	just,
universitet	university,
psykos	phychosis,
bollen	the ball,
viktigt	important,
human	human,
anders	anders,
beskriver	describes,
premiärminister	prime minister,
fysiker	physicist,
hävdar	assert,
bokstäver	letters,
troligt	likely,
hävdat	claimed,
självstyrande	independent,self-governance,
strax	soon,just,
julen	christmas,
jules	jules,
borgen	castle,the castle,
språkets	the language's,
arkitekturen	the architecture,
gustav	gustav,
särdrag	features,
följaktligen	consequently,
gustaf	gustaf,
trafikerar	frequent,
bekräftat	confirmed,
fastställdes	confirmed,
medborgarskap	citizenship,
kommunerna	the municipalities,
släkting	relative,
litauen	lithuania,
syrien	syria,
kemiska	chemical,
vattnet	the water,
kontinent	continent,
kunna	be able,
befolkningen	the population,
jupiter	jupiter,
befann	located,
kemiskt	chemically,
miljöproblem	environmental problem,environmental problems,
arthur	arthur,
däggdjuren	the mammals,
säsongerna	seasons,
shakespeare	shakespeare,
hertig	duke,
filmatiserats	cinematized,
benämns	is mentioned,
versionen	the version,
burj	burj,
versioner	versions,
bolt	bolt,
härstamma	stem,
burr	burr,
förkortat	shortened,
fördelen	the advantage,
därutöver	moreover,
omröstning	vote,
tolkats	interpreted,
tillverkas	manufacture,
strömmar	streams,flow,
grenen	the branch,
negativa	negative,
förknippade	associated,
äktenskap	marriage,
psykisk	psychic,
grundades	founded,was founded,
spåra	track,
havsnivån	sea level,
fastlandet	mainland,
märks	noted,
tennis	tennis,
könen	the sexes,
bönder	farmers,
bolivia	bolivia,
själv	alone,
byggnaden	building,the building,
berg	mountain,
japansk	japanese,
bero	depend,
epoken	the epoch,
sydligaste	southernmost,most southern,
spelade	played,
positiv	positive,
slaviska	slavic,
regeringen	the government,
båten	the boat,boat,
skelett	skeleton,
avsnitt	part,episode,
socialdemokrater	social democrats,
handelspartner	trading partner,
publiceringen	the publication,publishing,
vista	vista,
handen	hand,
handel	trade,
svärd	sword,
digital	digital,
kungamakten	the monarchy,
sades	was said,
överenskommelse	deal,
frodo	frodo,
exporten	the export,
accepterade	accepted,
rött	red,
riktad	directed,
ökande	increasing,
fss	fss,
expandera	expand,
riktat	pointed,
riktas	direct,
riktar	targets,
armar	arms,
bomben	the bomb,
telefon	telephone,
sanna	true,
manager	manager,
bomber	bombs,
vikingarna	the vikings,
dä	the elder,
imperiet	the empire,
avbrott	break,
uppdelning	partitioning,
petersburg	petersburg,
dö	die,
apartheid	apartheid,
trenden	the trend,
afrikansk	african,
höjdes	increased,was raised,
dit	there,
spets	point,
olympia	olympia,
ville	wanted,
malmö	malmö,
villa	house,villa,
reklamen	the commercial,
rymden	space,
utlösning	ejaculation,
hästen	the horse,
bakom	behind,
afghanistan	afghanistan,
viktig	important,
kokain	cocaine,
föredrog	preferred,
lönneberga	lönneberga,lonneberga,
somalia	somalia,
producent	producer,
tibet	tibet,
henry	henry,
köket	the kitchen,
avsaknad	absence,
beskrivits	described,
boy	boy,
diagnoser	diagnoses,
canadian	canadian,
bor	lives,
gyllene	golden,
folkmun	colloquially,
bok	book,
extrem	extreme,
mänsklighetens	humanity's,humanities,
diagnosen	diagnosis,the diagnose,
hotell	hotel,
sporter	sports,
utövar	exercise,
utövas	is practised,exercised,
världshälsoorganisationen	world health organization,
sporten	the sport,
religionsfrihet	religious freedom,
enormt	gigantic,
platån	sycamore,the plateau,
skräck	horror,
hemmaarena	home ground,
tennisspelare	tennis player,
semifinalen	semi finals,
kristian	kristian,
förbjöds	forbidden,
detaljer	details,
avsattes	dismissed,
brukade	used to,
kemisk	chemical,
fly	escape,
hände	happened,
tokyo	tokyo,
mästarna	the champions,
söka	search,
kombination	combination,
vittnen	witnesses,
akademien	academy,
präglade	characterized,
bristande	wanting,lack,
ulf	ulf,
hiroshima	hiroshima,
kenneth	kenneth,
uruguay	uruguay,
winston	winston,
agent	agent,
bemärkelse	meaning,
dennis	dennis,
oslo	oslo,
engelsmännen	the english,the british,
ekonomiska	economical,
till	to,
gitarrist	guitarist,
nye	new,
regeringstid	term of government,
överensstämmer	conform,
uppföljare	sequel,
läkare	doctor,
maj	may,
mao	mao,
man	one,
asien	asia,
sådana	such,
tala	speak,
block	block,
basket	basketball,
romantiken	romance,
sådant	such,
bevisa	prove,
alfabetet	the alphabet,
unionen	the union,
gällde	applied,
oktoberrevolutionen	october revolution,
moralisk	moral,
huvudsak	main thing,
motståndet	the resistance,the resistence,
verksam	active,
landskap	province,landscape,
sekter	sects,
äkta	genuine,
nazisterna	nazis,
växte	grew,
main	main,
texas	texas,
lägst	lowest,
steget	step,
janeiro	janeiro,
domstolar	courts,
vindkraft	wind power,
färg	colour,
uppskattning	appreciation,
tysklands	germanys,
hellre	rather,
vattendrag	streams,watercourse,
avkomma	offspring,
saudiarabien	saudi arabia,
canada	canada,
håkansson	hakansson,
pamela	pamela,
områdena	the areas,
tronföljare	successor,
kattdjur	felidae,cat,
ort	neighborhood,
konstnär	artist,
chiles	chile's,
dubbla	double,
snabbast	fastest,
miley	miley,
ord	word,
romarna	the romans,
anledning	reason,
självmord	self-killing,suicide,
rankningar	rankings,
dagsläget	present situation,
stängdes	closed,
centrala	central,
uttalanden	statements,
här	here,
rachel	rachel,
centralt	central,
skapandet	creation,the making,
kommunism	communism,
spänningen	exitement,
visas	shown,
västbanken	the west bank,
grundämnen	elements,
örebro	Örebro,
öronen	the ears,
besluten	decisions,
anus	ass,anus,
köpenhamns	copenhagen's,
fysiska	physical,
fysiskt	physical,
danny	danny,
löstes	solved,
drevs	was driven,
beslutet	the decision,
passade	suiting,suited,
fiender	enemies,
fienden	the enemy,
medlemmarna	the members,
lugn	calm,
fordon	vehicle,
marklund	marklund,
slöt	closed,
större	bigger,
tänder	teeth,
orsakerna	the causes,
kevin	kevin,
adeln	nobility,
nikola	nikola,
skulptur	sculpture,
centralbanken	central bank,
politiskt	political,
performance	uppträdande,
channel	channel,
norman	norman,
morden	murders,
politisk	political,
teoretiskt	theoretic,
ishockey	ice hockey,
civilisationer	civilizations,
otaliga	countless,
drottning	queen,
grammatik	grammar,
österut	eastwards,
kontrolleras	is controlled,
ungdom	youth,
civilisationen	civilization,
adolfs	adolf's,
generalsekreterare	secretary general,
helig	holy,
passande	fitting,suitable,matching,
historien	history,
statsmakten	the government,power,
medeltidens	medieval,
ges	be given,
ger	give,
klasser	classes,
kulturellt	cultural,
landets	the country's,
vintergatan	the milky way,
firade	celebrated,
rasen	the race,
himmlers	himmlers,
försörjning	sustentation,
bengtsson	bengtsson,
statistiska	statistical,
dianno	di'anno,dianno,
spridda	spread,
världskrigen	the world wars,
london	london,
tolfte	twelth,
relativt	relatively,
sekulära	secular,
fokuserar	focuses,
toppade	topped,
sean	seab,
stadsdelar	districts,city districts,
utgiven	published,
menar	means,
kandidater	candidates,
försvarsmakten	national defense,
personligt	personal,
personliga	personal,
august	august,
jr	junior,
åker	go,
timme	hour,
tum	inch,
lexikon	lexicon,
kirsten	kirsten,
rugby	american fotboll,
ån	the river,
tour	tour,
ås	ridge,
år	the year,year,
tryck	print,
vilja	will,
cancer	cancer,
statschefen	the head of state,
syntes	synthesis,
mätningar	measurements,measurments,
ryggen	the back,
barry	barry,
överföra	transfer,
mark	ground,
mars	march,
plötsligt	suddenly,
marx	marx,
mary	mary,
kultur	culture,
skriven	written,
cobain	cobain,
partido	partido,
avskaffa	abolish,
bmi	bmi,
spelfilmer	motion pictures,feature film,
skrivet	written,
fortsatt	continued,
dragit	dragged,
uppstod	developed,
kategorimän	category: men,
insåg	realized,
nionde	ninth,
intressanta	interesting,
uppmanade	urged,
liknande	similiar,similar,
sydkorea	south korea,
par	pair,
edwin	edwin,
lava	lava,
hålla	keep,
stött	met,
samt	also,as well as,
hösten	the fall,the autumn,
kuba	cuba,
teknisk	technical,
lösningar	solutions,
sömn	sleep,
wahlgren	wahlgren,
gates	gates,
bebyggelse	settlement,
dinosaurierna	dinasaurs,
skapelse	creation,
väst	west,the west,
byggnad	building,
reaktioner	reactions,
våld	violence,
jakten	the hunt,
ideologiskt	ideological,
bowie	bowie,
gotland	gotland,
ideologiska	ideological,
motverka	counteract,
trä	wood,
vintern	the winter,
mån	concerned,
mor	mother,
prägel	mark,
tillbehör	accessory,
jakt	hunt,
temperatur	temperature,
underarter	subspecies,
kollektiv	collective,
mod	courage,
adams	adams,
började	started,
födde	gave birth too,
manhattan	manhattan,
sågs	was observed,
göran	göran,
göras	be made,
feodala	feudal,
förr	sooner,
förs	led,
jordbruket	the agriculture,
fört	lead,
reportrar	reporters,
konsten	the art,
ända	as far as,
demokratisk	democratic,
samman	together,
moderata	moderate,
tunnlar	tunnels,
londons	london's,
cellen	the cell,
olof	olof,
akon	akon,
sjätte	sixth,
celler	cells,
allians	alliance,
metaforer	metaphores,
lands	on land,
lagarna	the laws,
retoriken	rhetoric,
newtons	newton's,
beskrivas	be described,
einstein	einstein,
intellektuella	intellectuals,
floderna	floods,
motivet	the motive,
behandling	treatment,
emellanåt	once in a while,
välmående	prosperous,
fullständiga	complete,
kvinnlig	female,
tillfälligt	temporarly,temporary,
eget	own,
utbredd	widespread,
egen	own,
vhs	vhs,
exemplar	example,
bibliografi	bibliography,
identifierade	identified,
parlament	parliament,
följde	followed,
youtube	youtube,
öns	the islands,
prestigefyllda	prestigious,
palats	palace,
sångerska	songstress,
goebbels	geobbels,
film	film,
genrer	genres,
effekt	effect,
spåren	the tracks,wake,
rubiks	rubik's,
vanligt	usual,
produktiv	productive,
stannade	stayed,
genren	genre,
faktorer	factors,
däremot	on the contrary,
ordna	arrange,
insats	stake,
ungarna	the young,
rykten	rumors,
ledning	guidance,
världsliga	worldly,
medicinska	medical,
palestinska	palestinian,
uppfostran	upbringing,
medicinskt	medical,
god	good,
snabbaste	fastest,
resolution	resolution,
åtskilda	separate,
mellanöstern	the middle east,
vila	rest,
hindrar	prevents,
liam	liam,
levern	the liver,
sund	sane,
symbolen	the symbol,
rwanda	rwanda,
symboler	symbols,
kasta	throw,
avhandling	thesis,
israeliska	isrealic,
stödja	support,
kulminerade	culminated,
miljoner	millions,
båtar	boats,
suttit	sat,
massor	lots,
publik	audience,
lärare	teacher,
värderingar	evaluations,
långhårig	long haired,
bebott	inhabited,
närhet	closeness,
jonas	jonas,
valt	chosen,
jackie	jackie,
tillkännagav	announced,
alexandria	alexandria,
sjukhuset	hospital,
varianterna	the diversities,
författaren	the author,
utmärkelsen	the award,
torra	dry,
diamond	diamond,
människa	man,
romersk	roman,
koma	coma,
tillkommer	reside,
hundraser	breed of dogs,
skivor	records,
vladimir	vladimir,
länkar	links,
roosevelt	roosevelt,
del	part,
baháulláh	bahullah,
samtliga	all,
hastigt	rapidly,fast,
latinets	the latin,
betoning	stress,
sjukdom	illness,
medförde	resulted,brought,
födseln	the birth,
sträng	string,
protein	protein,
makten	the power,
hämta	fetch,
psykotiska	psychotic,
stig	stig,
sammanfaller	coincides,
försvinner	disappears,
primära	primary,
vikten	importance,
makter	powers,
hoppade	jumped,
avtalet	the contract,
pettersson	pettersson,
laboratorium	laboratory,
huvudkontor	central office,headquarters,
vatten	water,
rastafarianer	rastafarian,
rockgrupper	rock bands,
paz	paz,
konservatismen	conservatism,
civila	civil,
inåt	inwards,
officiella	official,
fältet	the field,field,
göra	do,
baltikum	baltics,
officiellt	official,
människans	humans,mankinds,
längden	lenght,
diskussion	discussion,
wilhelm	wilhelm,
gustafsson	gustafsson,
suverän	terrific,
ställas	set,be set,
fängelse	prison,
sexuellt	sexual,
robbie	robbie,
kungarna	the kings,
namibia	namibia,
inleder	initiates,
anslöt	joined,
mental	mental,
fisk	fish,
flytta	move,
förenade	united,
energi	energy,
perry	perry,
sanningen	the truth,
östman	Östman,
oftast	most often,
infrastrukturen	infrastructure,
ölet	the beer,
forskning	research,
perro	perro,
fullständig	complete,
konflikt	conflict,
eventuellt	eventually,
investeringar	investments,
finland	finland,
styrs	ruled,
fått	was given,
styre	rule,
ensam	alone,
styra	steer,
säkerhetsråd	security council,
treenighetsläran	trinity,school of trinity,
snarast	rather,as soon as possible,
derivator	derivative,
kom	came,
lördagen	the saturday,
observationer	observations,
förhindrar	prevents,
park	park,
järnvägar	failways,
triangeln	the triangle,
gudarna	the gods,
domstolen	the court,
matteusevangeliet	gospel of matthew,
följden	result,
fort	quickly,
knapp	bare,
personens	the persons,
hellström	hellström,
baháí	bahá'í,
avtar	declines,
följdes	was followed,
försökte	tried,
gjord	made,
gjort	made,
mountain	mountain,
hundratals	hundreds of,hundreds,
infrastruktur	infrastructure,
caesar	caesar,
genast	immediately,
taktik	strategy,
lettland	latvia,
krafter	forces,
gillade	liked,
kraften	the force,
utbrott	outbreak,
laila	laila,
högt	high,
ko	cow,
km	kilometers,
kr	kronas,
liechtenstein	liechtenstein,
organisk	organic,
thomas	thomas,
venedig	venedig,
byttes	was exchanged,
relation	relation,
fina	beautiful,fine,
valet	the election,
antagit	presumed,
undre	lower,
wallenberg	wallenberg,
medverka	take part,participate,
tionde	tenth,
förbudet	the union,
avseende	regard,
blomstrade	flourished,
typiskt	typical,
notation	notation,
vänskap	friendship,
express	express,
förklarat	declare,
typiska	typical,
husen	the houses,
skickas	is sent,
skickar	sends,
brukar	usually,
boende	resident,
uttrycket	the expression,
uttrycker	expressing,
flykt	escape,
somrar	summers,
styrdes	governed,
suveränitet	sovereignty,
vind	wind,
godkännas	be approved,
landsbygden	rural area,
champagne	champagne,
romarriket	the roman empire,
bildandet	establishment,
framförs	is presented,
rörelserna	the movements,
kritiserades	critisized,
framföra	convey,
medlem	member,
musklerna	the muscles,
statligt	governmental,
uppfattning	understanding,
restaurang	restaurang,
romska	romani,
beta	graze,
globala	global,
kroatiens	croatias,
förklaring	explanation,
folkmord	genocide,
karaktären	character,
karaktärer	characters,
således	hence,thus,
tennessee	tennessee,
globalt	globally,
behöll	kept,
våningar	floors,
laos	laos,
bestämde	chose,
konspirationsteorier	conspiracy theories,
inför	before,
bengt	bengt,
popularitet	popularity,
gav	gave,
effektiva	effective,
gas	gas,
vana	familiar,
kalmar	kalmar,
effektivt	effective,
trupperna	troops,the troops,
detsamma	the same,
motorväg	highway,
åtalades	was prosecuted,
spridning	diffusion,distribution,
döptes	baptised,
portugal	portugal,
arenan	arena,
rederiet	the shipping company,shipping company,
dödar	kills,
dödas	killed,
administrationen	administration,
dödad	killed,
tyder	indicates,
sapiens	sapiens,
utmed	along,
skotska	scottish,
syd	south,
jerusalems	jerusalem's,
koloniala	colonial,
dopamin	dopamine,
nämnde	mentioned,
mot	against,
noll	zero,
kapitel	chapter,
albanien	albania,
jorderosion	earth erosion,
ministerrådet	minister counsellor,
norrland	norrland,
dikter	poems,
bibeln	bible,
passerar	passes,
alternativt	alternatively,alternative,
tropisk	tropical,
sparta	sparta,
administrativt	administrative,
monarkin	the monarchy,
administrativa	administrative,
åtal	prosecution,
dubbelt	double,
bil	car,
kejsaren	the emperor,
avlidna	diseased,
möttes	met,
bit	piece,
indonesiska	indonesian,
planeterna	the planets,
grå	grey,
kolonialtiden	the colonial times,
princip	principle,
möjlig	possible,
tillstånd	condition,
figurerna	characters,
google	google,
identisk	identical,
egyptiska	egyptian,
verkat	worked,
studerar	studies,
cocacola	coca cola,
västergötland	västergötland,
måste	have to,
per	per,
pratar	talks,talking,
självstyre	autonomy,self-governance,
energin	the energy,
lösningen	the solution,
därför	because,therefore,
ockuperade	occupied,
drama	drama,
fallit	fallen,
erkänner	admits,
styrelse	board of directors,
ontario	ontario,
turkiska	turkish,
medvetande	consciousness,
jaga	hunt,
serie	cartoon,
konsul	consul,
bostäder	residences,
jonathan	jonathan,
skillnaden	the difference,
ledningen	the lead,
planen	the plan,
planet	planet,
smycken	jewlery,
sultanen	sultan,
planer	plans,
frälsning	salvation,
reidar	reidar,
titel	title,
expedition	expidition,expedition,
förbjudna	forbidden,prohibited,
materia	materia,
tyskland	germany,
västerås	västerås,
voltaire	voltaire,
familjer	families,
årstiderna	the seasons,
familjen	the family,
makedonien	macedonia,
maos	mao's,
länders	countries',
samla	collect,
mutationer	mutations,
nådde	reached,
ritualer	rituals,
talades	spoken,spoke,
regionala	regional,
sambandet	the connection,connection,
dramatiker	dramatist,
judisk	jewish,
regionalt	regionally,
jason	jason,
stänga	close,
arvet	the inheritance,
penis	penis,
frankrike	france,
sigmund	sigmund,
stängt	closed,
intensivt	intensive,
privat	private,
medlemskap	membership,
sydafrikanska	south african,
sahlin	sahlin,
intensiva	intensive,
kollaps	collapse,
atlas	atlas,
graven	the grave,grave,
jakob	jakob,
luleå	luleå,
släppte	released,
tjänade	earned,
varnade	warned,
färöarna	the faroe islands,
beräkna	calculate,
exemplet	the example,
joel	joel,
reguljära	regular,
månens	the moon's,the moons,
warszawa	warsaw,
naturens	nature's,
joey	joey,
störtades	overthrown,
överhöghet	supremacy,
utbredda	widespread,
påsken	easter,
höjdpunkt	high point,
edison	edison,
går	goes,
chicago	chicago,
tillkomst	origin,
placering	placement,
vätet	the hydrogen,
och	and,
börja	start,
extrema	extreme,
mottagaren	the recipient,
populäraste	most popular,
sina	their,
honom	him,
svårigheter	difficulties,
skada	damage,
alaska	alaska,
katolicismen	catholisism,
lagförslag	bill,
miljard	billion,
färgade	colored,
protokoll	protocol,
uppnår	achieve,
uppnås	is achieved,
talare	spoke,
privata	private,
hennes	her,
nås	reached,
filippinerna	the philippines,
betraktar	regard,
nåd	mercy,grace,
lima	lima,
somrarna	summers,
kinesisk	chinese,
skotsk	scottish,
chi	chi,
gruppspelet	group play,
fånga	capture,
döpt	baptized,
söder	south,
geografisk	geographic,geographical,
titanics	titanic's,
iis	ii's,
prinsen	the prince,
ledamöterna	commisioners,
strider	battles,
utropade	cried out,
självständighet	independence,
iii	iii,
baserad	based,
baseras	based,based on,
baserat	based,
väldet	the rule,
indianerna	the indians,
titlar	titles,
mozarts	mozart's,
cecilia	cecilia,
fett	fat,
internationellt	internationally,
lanserade	introduced,
internationella	international,
rousseau	rousseau,
riktig	real,
klar	done,
billiga	cheap,
föddes	was born,
herrlandskamper	men's international contest,
mötte	met,
spannmål	grain,
klan	clan,
rådhus	courthouse,
billboardlistan	bilboardlist,
omslaget	the cover,
innebär	means,
industrier	industries,
la	la,
variationer	variations,
tvungna	forced,forced to,
weber	weber,
dag	day,
spektrum	spectra,
utfärdade	issued,
periodiska	periodic,
sammanhanget	context,
tolkade	interpreted,
day	day,
kontinuerligt	continuous,continous,
beslut	decision,
morris	morris,
syftade	alluded to,
lysande	brilliant,
krita	chalk,
humanism	humanism,
kristiansson	kristiansen,
dokumentär	documentary,
programmet	the application,
arbetskraft	workforce,labor,
nödvändiga	essential,
mats	mat's,
kärnan	core,
nödvändigt	neccessary,necessary,
deras	their,
återta	retake,
webbplats	website,
franz	franz,
odlas	cultured,
arbetare	workers,
längre	longer,
inleds	starts,
gravid	pregnant,
medelhavsområdet	the mediterranean region,the mediterranean area,
farbror	uncle,
fotografier	photographs,
nivå	level,
south	south,
liberaler	liberals,
stämmer	correct,
genomgår	undergoes,
uppger	states,
levnadsstandarden	the standard of living,
fruktade	feared,
omständigheter	circumstances,
veckan	the week,
utlopp	outflow,
energikällor	sources of energy,
drabbade	affected,
uppskattades	was appreciated,
leden	lines,the route,
demonstrationer	demonstrations,
bundna	tied,
stället	the place,
innehade	possessed,
firades	was celebrated,
sjögren	sjögren,
släkten	the family,
ställen	places,
bevarats	protected,
domaren	the judge,
matematisk	mathematical,
uteslutande	exclusivly,exclusively,
osmanska	osmanian,
mälaren	mälaren,
premiär	premiere,
aristoteles	aristoteles,
biologiska	biological,
älgar	moose,
följa	follow,
basist	bassist,
uganda	uganda,
idag	today,
följt	followed,
mil	swedish miles,
min	my,
skottland	scotland,
kroppar	bodies,
tidningar	magazines,
låg	low,
lån	loan,
konstverk	work of art,
konkurrerande	competing,
resurser	resources,
resultatet	the result,
dinosaurier	dinosaurs,
varandras	each others,
missionärer	missioners,
resultaten	the results,
sedan	since,
sist	last,
herman	herman,
republikanska	republican,
milano	milano,
deuterium	deuterium,
tidskrift	newspaper,
definiera	define,
styrka	power,
utgångspunkt	starting point,point of departure,
charles	charles,
inhemsk	native,
timmar	hours,
kurfursten	elector,
rumänska	romanian,
järnvägen	railroad,
euroområdet	eurozone,
rytmiska	rhythmic,
satan	satan,
organiska	organic,
snitt	on average,average,
arean	the area,
buddhismen	buddism,
uppehåll	hiatus,
richards	richards,
vinsten	the win,
organ	body,
nazitysklands	nazi germany,
majoriteten	the majority,
byggdes	was built,
national	national,
svenska	swedish,
egentlig	actual,
susan	susan,
seder	custom,
wembley	wembley,
bör	should,
terräng	terrain,
ordentligt	properly,
översikt	overview,
ronja	ronja,
industrialisering	industrialization,
uppskattade	estimated,appreciated,
stiga	rise,
hårdare	harder,
säkerheten	the security,
översättas	translated,be translated,
viktigare	more important,
hämtade	brought,
buddhas	buddhas,
konservativa	conservative,
miniatyr|karta	miniature|map,
återförening	reunion,
aktuellt	relevant,
kröntes	crowned,
aktuella	current,
kommendör	commandor,
fester	parties,
inneburit	meant,
befogenhet	warrant,authority,
tunisien	tunisia,
grupperingar	groups,
gaza	gaza,
asteroider	astroids,
försvar	defence,
stationen	station,
orange	orange,
västmakterna	western powers,
thåström	thastrom,
augusti	august,
bruket	the use,
stalin	stalin,
klassificera	classify,
dyker	dives,
tagits	taken,
fördrag	treaty,
partner	partner,
händelserna	the happenings,
lämnade	left,
blodtrycket	the blood pressure,
sångerna	the songs,
fler	more,
heinrich	heinrich,
hinduismen	hinduism,
kontrollera	control,
framförallt	above all,
kallas	called,
vanliga	regular,usual,
center	center,
öde	fate,
seth	seth,
sett	seen,
jupiters	jupiter's,
stores	the great's,
mystiska	mystical,
wagner	wagner,
grekiskans	greek,
flertal	majority group,
reformer	reformers,reforms,
mentala	mental,
landområden	land areas,
förnuft	reason,
uppmärksamhet	attention,
lika	similar,alike,
dubai	dubai,
koden	the code,
tusentals	thousands,
likt	like,
sarajevo	sarajevo,
works	works,
albumets	album's,
starkaste	the strongest,
profet	prophet,
etablerades	was established,
joachim	joachim,
skildras	is depicted,
definitionen	the definition,
definitioner	definitions,
starkare	stronger,
leopold	leopold,
about	about,
glada	happy,
tomt	empty,
andel	share,
värd	worth,
alexanders	alexanders,
förstärka	strengthen,
socken	parish,
omgiven	surrounded,
potatis	potato,
tränger	cut in,
skapade	created,
australiska	australian,
ljusare	lighter,
hatar	hate,
åter	again,
skog	wood,
kuben	the cube,
strävhårig	hispid,
föga	little,
förändrades	changed,
kväll	evening,
klockan	clock,o'clock,
brand	fire,
bröder	brothers,
kraft	power,
bud	bid,
vetenskap	science,
utrymme	space,
lissabon	lisbon,
australiens	australia's,
omfatta	cover,
kaffe	coffee,
minuter	minutes,
hästens	horses,
tolkningen	interpretetation,
omloppsbanor	orbits,
autism	autism,
kommuner	municipalities,
manlig	male,
proteiner	proteins,
uppfattar	percieves,
picchu	picchu,
stimulans	stimulating,
betonade	emphasized,
ljuset	the light,
försämrades	worsening,
astronomi	astronomy,
variation	diversity,
koncentrationsläger	concentration camp,
akademisk	academical,
philips	philips,
fakta	fact,
winnerbäck	winnerback,
baker	baker,
uggla	owl,
uppfattningen	comprehension,
framför	in front of,
förbundet	the union,
okänd	unknown,
slogs	fought,
påsk	easter,
antisemitiska	antisemetic,
anfallet	the attack,
paris	paris,
deltagit	participated,
kapacitet	capacity,
under	under,
nordost	the northeast,
ägande	owning,
jack	jack,
ovanstående	above,
minskat	decreased,has decreased,
öppna	open,
venus	venus,
verklig	real,
reklam	advertisement,
markerar	selects,
uppdelningen	division,
manus	script,
läget	location,
läger	camp,
stridigheter	oppositions,
drivande	driving,
ebba	ebba,
notera	note,
liberty	liberty,
aktiva	active,
zink	zinc,
språken	languages,
prata	talk,
medelhavsklimat	mediterranean climate,
beck	beck,
preparat	substance,
studio	studio,
atombomberna	the nuclear bombs,
sommartid	summer-time,during summer,
komplex	complex,komplex,
ty	for,
precis	precisely,
gällande	regarding,
koloniserades	is colonized,
upptäckter	discoveries,
upptäcktes	discovered,
julie	julie,
erektion	erection,
misslyckats	failed,
försvarsmakt	armed forces,
eftervärlden	the world,
mattias	mattias,
vinst	profit,win,
miniatyr|px|en	miniature,
konserterna	the concerts,
skicka	send,
behandlingar	treatments,
återstående	remaining,
muse	muse,
övertala	convince,persuade,
ludvig	ludvig,
ansökte	applied,
fermentering	fermentation,
rörelse	movement,
igelkottens	the hedgehog's,
henri	henri,
mm	millimeter,
arméns	the army's,
antiken	the ancient world,
mr	mr,
partiets	parties,
utlöste	triggered,
fröken	miss,
smält	melted,
väpnade	armed,
gata	street,
elektriskt	electric,
beskrev	depicted,described,
målen	goals,
förståelse	understanding,
mest	mostly,
västvärlden	western world,
målet	the target,
miniatyr|px|ett	miniature,
frågade	asked,
 cm	centimeters,
nagasaki	nagasaki,
kategorier	categories,
kubanska	cuban,
kontrollen	control,the control,
existera	exist,
arbetat	worked,
arbetar	work,works,
kejsare	emperor,
kampen	fight,
arresterades	was arrested,
vitt	widely,
besittningar	holdings,
frivillig	optional,
brinner	on fire,
edith	edith,
nytt	new,
blott	merely,
upptagen	occupied,
avskaffandet	abolishment,
jämförelser	comparison,
detroit	detroit,
sauron	sauron,
newport	newport,
storlek	size,
ursprungligen	originally,
platina	platinum,
nio	nine,
behövs	is needed,
kuwait	kuwait,
receptorer	receptors,
användningen	the use,
ammoniak	ammonia,
riktning	direction,
danmarks	denmark's,
paulus	paulus,
behöva	need,
independence	independence,
områdets	the area's,
kandidat	candidate,
fred	peace,
samlade	collected,
inom	within,
drygt	approximately,
statsministern	head of state,
studera	study,
tolerans	tolerance,
bredvid	next to,
vetenskapliga	scientific,
samhälle	society,
befolkade	populated,
vetenskapligt	scientifically,
transporterar	transports,
transporteras	is transported,
nyheter	news,
säsong	season,
museet	the museum,
föreslagits	was suggested,
nhl	nhl,
tillåts	is allowed,
återvände	returned,
sexuella	sexual,
×	x,
yngste	youngest,
punkten	point,
meddelanden	messages,
å	on,
ton	tone,
punkter	points,
tom	tom,
uppkommit	arisen,
tog	took,
adjektiv	adjective,
ifrågasatts	is questioned,
skildes	was seperated,
meddelande	message,
infaller	falls,
territoriella	territorial,
slutsats	conclusion,
mjölk	milk,
uppmuntrade	encouragement,encouraged,
nedgång	decline,fall,
rak	straight,
rör	touches,
störningar	disorder,
växer	grows,
ras	race,
motståndaren	the opponent,
industriellt	industrial,
hittats	found,
situationer	situations,
lanseringen	the release,
användning	use,
öarna	the islands,
industriella	industrial,
academy	academy,
situationen	situation,
mekaniska	mechanical,
tvingas	forced,
elektricitet	electricity,
fralagen	the fra law,
motsatt	opposite,
tanzania	tanzania,
sekt	sect,
metan	methane,
inflytande	influence,
flod	river,
utkanten	the outskirts,
idrott	sports,
järnvägarna	the railways,
queen	drottning,
gränserna	borders,
radio	radio,
earth	earth,
sagt	said,
radie	radius,
absolut	absolute,
turkar	turks,
claude	claude,
florens	florens,
vinna	win,
ägare	owner,
gods	domain,
holländska	dutch,
andras	others,
kommunisterna	the communists,
guatemala	guatemala,
gogh	gogh,
haiti	haiti,
ändras	be changed,
ursäkt	excuse,
ändrat	changed,
lovat	promised,
publicerades	published,
tidningen	the newspaper,
birgitta	birgitta,
kroppen	the body,
sakta	slowly,
ockuperat	occupied,
fördomar	prejudices,
kristendomen	chritianity,
antikens	ancient,
populär	popular,
slottet	the castle,
allra	most,
mun	mouth,
förhållande	in relation,
ordnade	arranged,
betonar	emphasize,
maniska	manic,
seden	the seed,
dödsorsaken	cause of death,
nummer	number,
kreativitet	creativity,
verka	operate,
misshandel	assault,
allierades	allied's,
begränsade	restricted,
förbränning	combustion,
avgöra	determine,
lägga	put,
grupper	groups,
solljus	sun light,
rumänien	romania,
reglera	expell,
möjliggjorde	allowed,
diktatorn	the dictator,
öster	east,
modernare	mor modern,
anspråk	claim,
spritt	spread,
invasionen	the invasion,
petrus	petrus,
depp	depp,
förståelsen	the understanding,
claes	claes,
nationer	nations,
därigenom	by which,thereby,
vojvodskap	voivodeship,
brott	crimes,
nationen	the nation,
kartan	the map,
äger	owns,
stadigt	steadily,
ökade	increased,
pekat	pointed,
negativ	negative,
welsh	welsh,
hundra	one hundred,
formatet	the format,
yngsta	youngest,
återvända	return,
gudom	deity,
dylan	dylan,
charlie	charlie,
spelad	played,
kemikalier	chemicals,
jean	jean,
spelat	played,
kraftigt	heavily,
järn	iron,
mängd	amount,
graden	rate,
europaparlamentet	the european parliament,
grader	degrees,
picasso	picasso,
utföras	performed,
kolväten	hydrocarbons,the hydrocarbon,
använt	used,
grundaren	the founder,founder,
aktiv	active,
regionerna	regions,
ekonomin	the economy,
tillgänglig	available,
auktoritet	authority,
uppträder	performs,
ladda	load,
modersmål	native language,
specifik	specific,
tillåtna	allowed,
fotbollen	soccer,
hund	dog,
gifter	marries,
lagstiftningen	law-making,
enat	united,
hushåll	household,
rådde	prevailed,
malaysia	malaysia,
besökt	visited,
motsatsen	the opposite,
ultraviolett	ultraviolet,
totalt	complete,wholly,
diktatur	dictator,
utse	name,
totala	total,
karaktäriseras	characterizes,
elitserien	elitserien,
monoteism	monotheism,
ishockeyspelare	ice hockey player,hockey players,
tillbringar	spends,
män	men,
spelare	player,
hotellet	the hotel,
meyer	meyer,
tvingades	forced,
systrar	sisters,
internationell	international,
tydliga	obvious,
primitiva	primitive,
civil	civil,civilian,
menade	meant,
systemet	the system,
tydligt	obvious,
isberg	ice berg,
sinne	mind,
lagt	laid,
kjell	kjell,
gia	gia,
metabolism	metabolism,
föreställa	imagine,
fadern	the father,
skulden	the guilt,
fängelsestraff	imprisonment,
italien	italy,
skulder	debts,
amerikanerna	the americans,
ruiner	ruins,
tillika	also,
araber	arabs,
regler	rules,
bildt	bildt,
hamn	harbor,
tronen	the throne,
judendomen	judaism,
förbud	ban,
liberalism	liberalism,
tätorten	conurbation,
tillverkade	manufactured,
ny	new,
tio	ten,
tid	time,
nr	number,
tätorter	conurbation,
nu	now,
phoenix	phoenix,
sätts	is placed,
tunna	thin,
kronprins	crown prince,
väckte	awakened,
beroendeframkallande	addictive,
rom	rome,
ron	ron,
rod	rod,
dvärg	dwarf,
knutsson	knutsson,
koreanska	korean,
udda	odd,
laura	laura,
mottagarens	the reciever,the receivers,
konstitutionell	constitutional,
federation	federation,
varvid	in which,
underhållning	entertainment,
flytt	escaped,
krossa	crush,
metod	method,
brother	brother,
olyckor	accidents,
beräknades	estimated,
tillverkningen	production,the production,
heinz	heinz,
trend	trend,
stilar	styles,
svartån	svartån,
förorter	suburbs,
port	gate,
ifråga	with regards to,
sociala	social,
månaderna	months,
angelina	angelina,
gräs	grass,
kamp	fight,
vindkraftverk	wind turbine,
enkla	simple,
metaller	metals,
angående	concerning,
turister	tourists,
lokal	local,
ankomst	arrival,
filmen	the movie,
tilltagande	increasing,
etablera	establish,
trummor	drums,
bolaget	the company,
russell	russell,
ande	spirit,
inblandade	involved,
kurder	kurds,
australian	australian,
turné	tour,
veckorna	weeks,
typerna	the types,
kär	in love,
övergå	transition,transend,
piano	piano,
styras	steered,
drabbades	affected,
läkemedel	medicine,
partnern	the partner,
rådgivare	counsellor,
valla	valla,
allvarlig	serious,
domkyrka	cathedral,abbey,
generell	general,
musikaliskt	musical,
springsteens	springsteens,
uppväxt	growing up,
bönorna	beans,
utdelades	distributed,
hemligt	secret,
hemliga	secret,
lätta	lighten,
avrättning	execution,
frivilliga	volunteers,
stöter	thrust,
simning	swimming,
muslimerna	the muslims,
inriktad	intent,
tvserien	the tv show,television program,
fascism	fascism,
sydliga	southern,
familjens	the familys,
flög	flew,
fenomen	phenomenon,
leva	live,
utrikespolitiska	foreign policy,
olika	different,
marknad	market,
persons	persons,
komplicerad	complicated,
orter	locations,
kartor	maps,
orten	the suburb,
komplicerat	complicated,
böcker	books,
utvecklingen	the development,
organisation	organization,
behandlingen	the treatment,the treament,
försvaret	the defense,
marleys	marley's,
hergé	herge,
femte	fifth,
hamilton	hamilton,
tredjedel	a third,
hotar	threatens,
opera	opera,
namn	name,
futharkens	the futhark's,
viggo	viggo,
hotad	threatened,
färger	colors,
bildning	education,form,
semifinal	semi finals,
stående	standing,
amerikansk	american,
behandlar	treat,
behandlas	treated,
upprepade	repeated,
stortorget	stortorget,
årliga	annual,
profil	profile,
accepterar	accepts,
accepterat	accepted,
kent	kent,
variant	variant,variety,
juldagen	christmas day,
zuckerberg	zuckerberg,
nått	reached,
hjalmar	hjalmar,
gallien	gaul,
produktionen	the production,
arbetet	the work,
traditionen	the tradition,
traditioner	traditions,
place	place,
politiken	the politics,
arbeten	works,
origin	origin,
begår	commits,
såldes	sold,
kontrollerade	controlled,
vågor	waves,
okända	unknown,
bahamas	bahamas,
givet	granted,
personlighetsstörningar	personality disorders,
spelats	been played,played,
kronprinsessan	crown princess,
montenegro	montenegro,
kallade	called,
hur	cage,
hus	house,
population	population,
smeknamn	nickname,
modellen	the model,
marinen	navy,marines,
löfte	promise,
kontroll	control,
framställning	production,
övertogs	overtaken,
modeller	models,
bildades	was formed,
hjärtat	the heart,
afrikanska	african,
anc	anc,
kromosomerna	the chromosomes,
maten	the food,
jordskorpan	earth crust,
världen	the world,
avstånd	distance,
förste	the first,
förhållandena	conditions,the conditions,
gustavs	gustavs,
konsert	concert,
stjärnornas	the star's,
knutna	associated,tied,
diskussioner	discussions,
falla	fall,
fria	free,
täcks	covers,
lisbet	lisbet,
elektromagnetisk	electromagnetic,
stövare	hound,
herren	the lord,
ronaldinho	ronaldinho,
mänskligheten	humanity,
sjunka	descend,
tror	believe,
bandets	the bands,
berättelsen	the story,
guld	gold,
flydde	fled,
ovanligt	unusual,
iväg	away,
ovanliga	unusual,
larsson	larsson,
jazz	jazz,
ansågs	seemed,
beredd	prepared,
tränade	trained,
dramat	the drama,
joker	joker,
republika	republic,
osäkert	insecure,uncertain,
förmån	benefit,
minnen	memories,
underlätta	ease,
stanley	stanley,
freden	the peace,
fredspriset	peace prize,peace price,
skett	happened,
önskade	wished,
återigen	yet again,
hämtat	collected,taken,
konstnären	the artist,
bekämpa	fight,
dödade	killed,
sydeuropa	southern europe,
region	region,
ordagrant	literal,
spindlar	spiders,
lenins	lenin's,
gjorde	did,
gjorda	made,
pakistan	pakistan,
utgåvor	issues,
period	period,
pop	pop,
fransk	french,
werner	werner,
statens	the government's,
utformning	layout,
hävda	claim,
poe	poe,
skånska	scanian dialect,scanian,
folken	the peoples,
strikta	strict,
förekomsten	existence,presence,
dagarna	the days,
musikstil	music style,
folket	the people,
invaderade	invaded,
anderna	the andes,
andres	andres,
andrew	andrew,
kapitulation	surrender,capitulation,
minister	minister,
använder	uses,
användes	was used,
cash	cash,
arnold	arnold,
spreds	spread,
fiende	enemy,
grundlagen	the constitutional law,
pippi	pippi,
kuriosa	trivia,
theta	theta,
knyta	tie,
grönland	greenland,
status	status,
fysiologi	physiology,
protoner	protons,
hjärta	heart,
linjerna	the lines,
göring	goring,
privilegier	privileges,
relaterade	related,
medvetna	aware,
kommunistisk	communistic,communist,
breda	wide,
without	without,
medellivslängd	average lifespan,life expectancy,
möta	meet,
helsingfors	helsingfors,
listorna	the lists,
kommentarer	comments,
förklarades	was explained,
allmän	general,
möte	meeting,
harrison	harrison,
moçambique	mozambique,
leta	search,
utvinns	extracted,
tim	tim,h,
rose	rose,
regent	regent,
rosa	pink,
utbyte	trade,
feminism	feminism,
vampyren	the vampire,
delhi	delhi,
utrikespolitik	foreign affairs,
möts	meets,
vampyrer	vampires,
riken	the kingdoms,
kommentar	comment,
afrikas	africas,
patrick	patrick,
anföll	attacked,
rammstein	rammstein,
styrkor	strenghts,
teorin	the theory,
gång	time,
passera	pass,
latinet	latin,
alkoholer	alcohols,
verksamheter	operations,businesses,
försvarare	defender,
tiders	days',
sitta	sit,
stopp	stop,
lärda	savants,
buddha	buddha,
antika	ancient,
uppbyggnad	construction,
willy	willy,
geografi	geography,
tyskt	german,
tyske	german,
on	on,
om	if,
indianska	native american,
spelet	the game,
of	av,
oc	oc,
stand	stand,
os	os,
spelen	the games,
befäl	command,
koppling	connection,
cambridge	cambridge,
beskrivning	description,
burton	burton,
trådlös	wireless,
medlemsstaternas	member state,
valley	valley,
genomfört	carried out,
jul	christmas,
inriktning	direction,orientation,
ekonomi	economy,
poes	poe's,
chaplin	chaplin,
kvinnornas	womens,
felix	felix,
närmast	closest,
fjorton	fourteen,
pontus	pontus,
operation	operation,
köpenhamn	copenhagen,
många	many,
utgifter	expenses,
babylon	babylon,
visade	showed,
grupp	group,
ockupation	occupation,
symbol	symbol,
erövring	conquest,
missbruk	abuse,
calle	calle,
visby	visby,
ali	ali,
alf	alf,
separat	seperate,separate,
ale	ale,
stödde	supported,
samhällen	communities,societies,
sakrament	sacrament,
gärning	deed,
funktionerna	the functions,
röstade	voted,
påstående	assumption,
kvar	left,
löper	runs,
oavgjort	draw,
far	father,
fas	phase,
runtom	throughout,around,
simpsons	simpsons,
sony	sony,
unionens	the union's,
tjeckiska	czech,
list	cunning,
kopplas	connected,
förtryck	opression,
lisa	lisa,
grekland	greece,
ted	ted,
istiden	the ice age,
tex	for example,
haag	the hague,
what	what,
spelning	gig,
upptäcka	discover,
regerade	reigned,
leeds	leeds,
upptäckt	discovered,discovery,
norden	the nordic countries,
soloalbum	solo album,
kärnvapen	nuclear weapons,
tillhörde	belonged to,
magnitud	magnitude,
arabemiraten	united arab emirates,
påföljande	subsequent,
filmerna	the movies,
stöd	support,
dahlén	dahlén,
syfta	aim,
socialdemokraterna	members of the social democracy,
anarkism	anarchism,
fängslade	imprisoned,
branden	the fire,
förebild	role model,
autonom	independent,
gemensamt	in common,
israel	israel,
permanenta	permanent,
cellerna	the cells,
akademiens	the academy's,
floyd	floyd,
östra	eastern,
naturligt	natural,
legender	legends,
salvador	salvador,
decenniet	decade,
kryddor	spices,
naturliga	natural,
duett	duet,
bosatt	resident,lived,
historiskt	historic,historical,
breaking	breaking,
brittisk	british,
satanism	satanism,
härstamning	origin,descent,
rocksångare	rock singer,
böhmen	bohemia,
grundämne	element,
fötterna	feet,
fötts	born,borned,
regnar	rains,
anarkistiska	anarchist,
praktiska	practical,
tsar	tsar,
homosexuella	homosexual,
grande	grand,
människors	humans,
instabil	unstable,
september	september,
gudarnas	the gods',
australien	australia,
längd	length,
lyder	obeys,
handlar	concerns,
abbey	abbey,
rikt	rich,
prag	prague,
stephen	stephen,
argentina	argentina,
fenomenet	the phenomenon,
dickens	dicken's,
medborgerliga	civil,
kärna	core,
postumt	posthumously,
marcus	marcus,
försöken	the tries,
journalisten	the journalist,
journalister	journalists,
försöker	tries,trying,
tvister	disputes,
ringar	rings,
betyg	grades,
sätt	way,
stenar	stones,
ollonet	the glans,
därvid	therewith,
väg	way,
vän	friend,
poliser	police,
ökad	increase,increased,
ersatt	replaced,
ökat	increased,
trummisen	the drummer,
fallet	the case,
stavningen	the spelling,
konsumtionen	consumption,
fallen	cases,
aminosyror	amino acids,
pablo	pablo,
bland	including,
blanc	blanc,
story	story,
misslyckas	fails,
stort	big,
motiveringen	the motivation,
storm	storm,
kristendomens	christianity's,
brasiliens	brazil's,
ecuador	ecuador,
mikael	mikael,
gränser	borders,
hotel	hotel,
kongress	congress,
serotonin	serotonin,
framtiden	the future,
fattigaste	the poorest,
gränsen	border,
siffra	number,
illegala	illegal,
matcherna	the games,
direkt	direct,
kina	china,
guden	the god,
stjärnan	the star,
kategorin	the category,
klubb	club,
anläggningar	facilities,
kusin	cousin,
tilldelas	assigned,
omskärelse	circumcision,
slåss	fight,
 km	kilometers,
bedriver	operate,
unga	young,
jämförelsevis	in comparison,
judas	judas,
judar	jews,
folkgrupper	ethnic groups,
electric	electic,
dagliga	daily,
stjärnans	the stars,
dagligt	daily,
industrialiserade	industrialized,
sånger	songs,
mineral	mineral,
influensan	the influenza,
sången	the song,
statsskick	polity,
kosovo	kosovo,
ursprungliga	original,
kolonialism	colonialism,
tilly	tilly,
månen	the moon,
tills	until,
beräkningar	calculations,
hit	to here,here,
hiv	hiv,
inklusive	including,
vardera	each,
händer	hands,
himmler	himmler,
solsystemet	the solar system,
utvidgade	expanded,
tvkanaler	tv channels,
mediciner	medicines,
avtal	contract,
tidszon	timezone,time zone,
vincent	vincent,
norrköping	norrköping,
virginia	virginia,
utsatt	exposed,
etiopien	ethiopia,
art	kind,
bart	bart,
fiske	fishing,
arg	angry,
arm	arm,
pär	pär,
planeras	is planned,
överföring	transfer,
uppskatta	appreciate,
inga	no,
planerat	planned,
planerad	planned,
latin	latin,
verksamhet	work,
där	where,
intäkter	incomes,
herrar	men,
uppkom	arose,
tiderna	the times,
startades	started,
lyssnar	listen,
hypotesen	the hypothesis,
lära	get to know,
sweet	söt,
vidare	moreover,
lärt	learned,
stärktes	was strenghten,
belägna	located,
östtyskland	east germany,
hypoteser	hypothesis,
ps	ps,
java	java,
skrev	said,
kungafamiljen	the royal family,
johannes	johannes,
inkluderas	is included,
byxor	pants,
resultat	result,results,
pi	pi,
chandler	chandler,
flight	flight,
togs	taken,
sydafrikas	south africa's,
rättigheterna	the rights,
konflikter	conflicts,
deltog	participated,
inspelningar	recordings,
ris	rice,
sjöarna	the lakes,
byggnaderna	the buildings,
skeppen	the ships,
fysisk	physical,
demografi	demographics,
tidpunkten	the time,the moment,
ideologier	ideologies,
listor	lists,
förföljelse	persecution,
spears	spears,
bröllopet	the wedding,
byar	villages,
uppbyggd	built-up,
författare	author,
sökte	searched,
kokpunkt	boiling point,
visats	shown,
italiensk	italian,
sjunga	sing,
vetenskapen	the science,
kyrkans	the church's,
uttalande	statement,
komplett	complete,
konstitution	constitution,
press	press,
remmer	remmer,
prince	prince,
skalv	quake,
minoriteter	minorities,
bostad	lodge,
omedelbar	immediate,
skall	shall,
minoriteten	minority,
emigrerade	emigrated,
synnerhet	specially,particular,
djupare	deeper,
begravdes	buried,
användas	used,
stoppade	stopped,
upplevelse	experience,
exakt	accurately,
våldsamma	violent,
näringsliv	business,
hittades	was found,
hittas	found,
minskning	decline,
norrut	north,
sjöfart	sea voyage,
kongo	congo,
trummis	drummer,
krigare	warrior,
låtarna	the songs,
föräldrar	parents,
grekerna	greek,
statyn	the statue,
anne	anne,
trinidad	trinidad,
anna	anna,
höjder	altitudes,heights,
turism	tourism,
palmes	plame's,
ställningen	position,
presenteras	presented,
judendom	judaism,
kostnaderna	the costs,
grundläggande	primary,
finansieras	financed,
tätt	tightly,
utropades	proclaimed,
dialog	dialogue,
täta	close,
socialistisk	socialistic,
sällsynta	rare,
medborgarna	the citizens,
hållet	way,
abbas	abbas,
km²	square kilometre,
håller	holds,
uppvisar	shows,
fast	even though,
jugoslavien	yugoslavia,
bruk	use,
organiserade	organized,
regionen	the region,
kombinationer	combinations,
sköter	handles,
regioner	regions,
junior	junior,
karolinska	caroline,
planeternas	the planets,planets,the planets',
angels	angels,
styrande	rulers,
erövrades	concoured,
guyana	guyana (name),
tolka	interpret,
z	z,
tidens	time's,
svenskspråkiga	swedish speaking,
tidpunkt	date,
däribland	including,
stadion	stadium,
psykoterapi	psychotherapy,
använts	was used,
mötet	the meeting,
möter	meets,
skyddar	protects,
sutra	sutra,
beräknar	values,
tittarna	the viewers,
medina	medina,
konvertera	convert,
råkar	happens to,
kaspiska	caspian,
oväntat	unexpected,
vice	vice,
europeiska	european,
nasa	nasa,
lagstiftning	law-making,
nash	nash,
steve	steve,
jimi	jimi,
stieg	stieg,
kolonialismen	the colonialism,
simon	simon,
uppmaning	exhortation,
fortfarande	still,
romerna	the romani,the romani people,
generella	general,
hinduism	hinduism,
fotnoter	footnotes,
varierar	varies,
vapen	weapon,
georgien	georgia,
medverkade	participated,
kommitté	committee,
avslutas	close,ends,
avslutat	completed,
historikern	historian,
byggt	built,
noter	notes,
utanför	outside,
musikaliska	musical,
melodier	melodies,
demokratiska	democratic,
bygga	build,
åtta	eight,
influerad	influenced,
anderssons	anderssons,
århundraden	centuries,
västlig	western,
konstant	constant,
folk	people,
influerat	influenced,
hölls	was held,
assisterande	assisted,
skrivna	written,
judy	judy,
dramatiska	dramatic,
bröts	was fractured,
koloni	colony,
hdmi	hdmi,
producenten	the producer,
diamanter	diamonds,
åtgärder	measures,
filosofi	philosophy,
astrid	astrid,
tvingats	forced,
buddhistiska	buddhistic,
ukraina	ukraine,
metro	metro,
innehar	holds,
elektronik	electronics,
anpassat	adapted,
plattan	plate,
översättningar	translations,
tjänar	earns,
zlatan	zlatan,
gemenskap	fellowship,
motor	engine,
varpå	whereupon,
from	from,
bestämmelser	measures,
usa	usa,
fel	errors,
fem	five,
sevärdheter	attractions,
inlandet	inland,
sorg	grief,
uran	uranium,
införande	introduction,
hindrade	prevented,
vägrade	refused,
slutade	quit,
beskriva	describe,
automatiskt	automatic,
tar	takes,
tas	is taken,
föreslår	suggest,
platser	places,
crick	crick,
platsen	place,
tag	while,
kanadensiska	canadian,
sir	sir,
ondska	evil,
beyoncé	beyoncé,
brian	brian,
undantaget	except,
sin	its,
väpnad	armed,
oavsett	regardless,
tack	thanks,
religiös	religious,
bertil	bertil,
frivilligt	voluntarily,
kontroversiella	controversial,
eritrea	eritrea,
light	light,
kommunikationer	communications,
besegrat	defeated,
skapande	creative,
elin	elin,
karlstad	karlstad,
blandas	mixes,
spotify	spotify,
listan	the list,
uppmärksammad	noticed,
floder	rivers,
permanent	permanent,
genomsnittlig	average,
lärjungar	disciple,
uppmärksammat	noticed,
cypern	cyprus,
betalade	payed,paid,
underjordiska	underground,
material	material,
östtimor	east timor,
växande	growing,
studios	the studio's,
wallander	wallander,
säsonger	seasons,
byter	changes,exchanges,
kvarteret	the neighborhood,
säsongen	season,
arterna	the species,
kritik	criticism,critisism,
förbjuda	ban,
svag	weak,
minskad	decreased,
hantverkare	craftsman,handy worker,
svar	response,
tagit	taken,
plural	plural,
förutsättningar	prerequisites,condition,
hörs	heard,
hört	heared,
vulkanutbrott	vulcano eruption,
lösas	solved,
york	york,
van	van,
philip	philip,
domare	judge,
hörn	corner,
fotbollslandslag	national football team,
gångna	past,
tyst	quiet,
barns	childrens,
via	through,
adrian	adrian,
tvserier	tv shows,
rudolf	rudolf,
ovanpå	on top of,
revolutionens	the revolutions,
isbn	isbn,
brasilien	brazil,
nietzsches	nietzsche's,
mått	measurement,
skyddade	protected,
nätverk	network,
åtskilliga	several,
fågelhundar	bird dogs,
förkortning	abbreviation,
merkurius	mercury,
omfattning	extent,
sankta	sankta,
rösträtt	right to vote,
valde	chose,
valda	chosen,
vingar	wings,
juli	july,
väntan	awaiting,waiting,wait,
dödligheten	mortality,
resterande	remaining,
holland	holland,
franske	the french,
utvisning	penalty,
framgång	success,
algeriet	algeria,
franskt	french,
tomma	empty,
tyskarna	the germans,
farliga	dangerous,
flyttat	moved,
cohen	cohen,
benny	benny,
avgörs	decided,is determined,
blir	become,
gäng	group,
intervju	interview,
byggas	build,
uppfann	invented,
lopp	race,
ansåg	thought,considered,
besittning	dominion,
protesterade	protested,
centra	center,
centre	centre,
who	who,
landslaget	the national team,
intogs	was captured,
staternas	states,
öken	desert,
planerade	planned,
förbundsrepubliken	the federal republic,
undersökte	investigated,
regeringschef	government,
miljontals	millions,
generna	the genes,
moberg	moberg,
blandade	mixed,
debatt	debate,
pastoral	pastoral,
eiffeltornet	the eiffel tower,
dödades	were killed,
asterix	asterix,
filmer	movies,
beroende	dependent,
allmänhet	in general,general,
träffa	meet,
gudar	gods,
presley	presley,
närstående	relative,kindred,
städer	cities,
begäran	request,
förbinder	connects,
mestadels	mostly,
nationernas	the nations,
motståndare	opponents,
anlände	arrived,
funktion	function,
betydande	important,
praktisk	practical,
vandrar	wanders,
joe	joe,
jon	jon,
barrett	barett,
influenser	influences,
påtagligt	substantially,
västerländsk	western,
brons	bronze,
vattnets	the water's,the waters,
bronx	the bronx,
förespråkare	spokesman,
betecknar	denotes,
betecknas	denote,
demens	dementia,
vittne	witness,
publicerad	published,
walt	walt,
innebära	mean,
framträdanden	appearances,
publicerat	published,
demografiska	demographic,demographical,
dödshjälp	euthanasy,
kopplade	connected,
mångfald	variety,
månar	moons,
marilyn	marilyn,
klart	done,
månad	month,
strindbergs	strindberg's,
naturtillgångar	natural resources,
pengar	money,
nickel	nickel,
klassen	the class,
turneringen	the tournament,
försvann	disappeared,
fortsättningen	the continuation,
plikter	duties,
godkännande	approval,
bråk	fights,
officiell	official,
största	biggest,largest,
anpassa	adjust,
fördelade	divided,
wild	wild,
explosionen	the explosion,
bekräftade	confirmed,
syftar	refers,seek to,
motiv	motif,
jehovas	jehovas,jehova's,
röra	move,
uppstå	develop,
ramels	ramel's,
buddhism	buddhism,
pojkar	boys,
samband	connection,
odlade	grew,
skickade	sent,
annekterade	annexed,
kustlinje	coastline,
övervägande	predominant,
romeo	romeo,
romer	romani people,
student	student,
misstag	mistake,
klubbar	clubs,
vilar	rests,
banden	the bound,
närma	approach,
ekosystem	ecosystem,
organisationens	the organizations,
rachels	rachel's,
erfarenheter	experience,
högskolor	colleges,
förtroende	confidence,
miljöer	environments,
antisemitism	antisemitism,
rocken	rock,
brutit	broken,
mytologiska	mythological,
jarl	jarl,
genombrottet	breakthrough,
alldeles	completely,
hoppa	drop out,
sky	sky,
rättsliga	legal,
engelsk	english,
ske	happen,
ska	will,
fyller	turns,
sanskrit	sanskrit,
färgen	the color,
älska	love,
nathan	nathan,
budet	the bid,the commandment,
miami	miami,
djupa	deep,
huruvida	whether,
sälja	sell,
påtryckningar	pressures,
säkra	reliable,safe,
juni	june,
tjeckoslovakien	czechoslovakia,
bibliska	biblican,
gäst	guest,
export	export,
högst	highest,
planering	planning,
gammalt	old,
setts	seen,
låter	let,
låten	the song,
sjunker	sinks,
äta	eat,
utsöndras	exudes,
uppvärmning	heating,warming,
mitt	my,
slut	end,
sommarspelen	summer games,
ljung	heather,
låna	borrow,
upplöstes	dissolved,
substantiv	noun,
tillräcklig	sufficient,enough,
överlevde	survived,
bestämma	decide,
greve	earl,
saken	the thing,
saker	things,
främre	front,
egna	own,
återvänt	returned,
någorlunda	fairly,
tillbringade	spent,
mäts	is measured,
en	a,
floden	the river,
vidta	take,
konstruktion	construction,
födelsetal	birthrate,birth rate,
val	choice,
upprättas	establish,
mäter	measuring,
nordamerikanska	north american,
lundell	lundell,
hundratal	hundred,
ingått	entered,
nödvändigtvis	by necessity,necessarily,
karta	map,
rybak	rybak,
tema	theme,
missnöjet	grievance,
inledning	introduction,
jenny	jenny,
reaktorn	reactor,
problemet	the problem,
stormakter	world powers,
utöva	exercise,
resultera	result,
illinois	illinois,
book	book,
ursprunget	origin,
åren	the years,years,
intresse	interest,
serbiska	serbian,
tolkas	is interpreted,interpret,
tolkar	interprets,
personligen	personally,
ställningar	positions,
markant	considerably,
stadens	the town's,the citys,
spontant	spontaneous,
bysantinska	byzantine,
tidning	newspaper,
